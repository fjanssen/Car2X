// nios_system.v

// Generated using ACDS version 12.1 177 at 2014.06.16.15:30:22

`timescale 1 ps / 1 ps
module nios_system (
		output wire [11:0] sdram_communication_wire_addr,                    //                  sdram_communication_wire.addr
		output wire [1:0]  sdram_communication_wire_ba,                      //                                          .ba
		output wire        sdram_communication_wire_cas_n,                   //                                          .cas_n
		output wire        sdram_communication_wire_cke,                     //                                          .cke
		output wire        sdram_communication_wire_cs_n,                    //                                          .cs_n
		inout  wire [31:0] sdram_communication_wire_dq,                      //                                          .dq
		output wire [3:0]  sdram_communication_wire_dqm,                     //                                          .dqm
		output wire        sdram_communication_wire_ras_n,                   //                                          .ras_n
		output wire        sdram_communication_wire_we_n,                    //                                          .we_n
		output wire [7:0]  pio_communication_led_external_connection_export, // pio_communication_led_external_connection.export
		input  wire        reset_reset_n,                                    //                                     reset.reset_n
		input  wire        clk_clk,                                          //                                       clk.clk
		input  wire [3:0]  tse_mac_conduit_connection_rgmii_in,              //                tse_mac_conduit_connection.rgmii_in
		output wire [3:0]  tse_mac_conduit_connection_rgmii_out,             //                                          .rgmii_out
		input  wire        tse_mac_conduit_connection_rx_control,            //                                          .rx_control
		output wire        tse_mac_conduit_connection_tx_control,            //                                          .tx_control
		input  wire        tse_mac_conduit_connection_tx_clk,                //                                          .tx_clk
		input  wire        tse_mac_conduit_connection_rx_clk,                //                                          .rx_clk
		input  wire        tse_mac_conduit_connection_set_10,                //                                          .set_10
		input  wire        tse_mac_conduit_connection_set_1000,              //                                          .set_1000
		output wire        tse_mac_conduit_connection_ena_10,                //                                          .ena_10
		output wire        tse_mac_conduit_connection_eth_mode,              //                                          .eth_mode
		output wire        tse_mac_conduit_connection_mdio_out,              //                                          .mdio_out
		output wire        tse_mac_conduit_connection_mdio_oen,              //                                          .mdio_oen
		input  wire        tse_mac_conduit_connection_mdio_in,               //                                          .mdio_in
		output wire        tse_mac_conduit_connection_mdc                    //                                          .mdc
	);

	wire          tse_mac_receive_endofpacket;                                                                                    // tse_mac:ff_rx_eop -> sgdma_rx:in_endofpacket
	wire          tse_mac_receive_valid;                                                                                          // tse_mac:ff_rx_dval -> sgdma_rx:in_valid
	wire          tse_mac_receive_startofpacket;                                                                                  // tse_mac:ff_rx_sop -> sgdma_rx:in_startofpacket
	wire    [5:0] tse_mac_receive_error;                                                                                          // tse_mac:rx_err -> sgdma_rx:in_error
	wire    [1:0] tse_mac_receive_empty;                                                                                          // tse_mac:ff_rx_mod -> sgdma_rx:in_empty
	wire   [31:0] tse_mac_receive_data;                                                                                           // tse_mac:ff_rx_data -> sgdma_rx:in_data
	wire          tse_mac_receive_ready;                                                                                          // sgdma_rx:in_ready -> tse_mac:ff_rx_rdy
	wire          sgdma_tx_out_endofpacket;                                                                                       // sgdma_tx:out_endofpacket -> tse_mac:ff_tx_eop
	wire          sgdma_tx_out_valid;                                                                                             // sgdma_tx:out_valid -> tse_mac:ff_tx_wren
	wire          sgdma_tx_out_startofpacket;                                                                                     // sgdma_tx:out_startofpacket -> tse_mac:ff_tx_sop
	wire          sgdma_tx_out_error;                                                                                             // sgdma_tx:out_error -> tse_mac:ff_tx_err
	wire    [1:0] sgdma_tx_out_empty;                                                                                             // sgdma_tx:out_empty -> tse_mac:ff_tx_mod
	wire   [31:0] sgdma_tx_out_data;                                                                                              // sgdma_tx:out_data -> tse_mac:ff_tx_data
	wire          sgdma_tx_out_ready;                                                                                             // tse_mac:ff_tx_rdy -> sgdma_tx:out_ready
	wire          nios2_communication_instruction_master_waitrequest;                                                             // nios2_communication_instruction_master_translator:av_waitrequest -> nios2_communication:i_waitrequest
	wire   [27:0] nios2_communication_instruction_master_address;                                                                 // nios2_communication:i_address -> nios2_communication_instruction_master_translator:av_address
	wire          nios2_communication_instruction_master_read;                                                                    // nios2_communication:i_read -> nios2_communication_instruction_master_translator:av_read
	wire   [31:0] nios2_communication_instruction_master_readdata;                                                                // nios2_communication_instruction_master_translator:av_readdata -> nios2_communication:i_readdata
	wire          nios2_communication_instruction_master_readdatavalid;                                                           // nios2_communication_instruction_master_translator:av_readdatavalid -> nios2_communication:i_readdatavalid
	wire          nios2_communication_data_master_waitrequest;                                                                    // nios2_communication_data_master_translator:av_waitrequest -> nios2_communication:d_waitrequest
	wire   [31:0] nios2_communication_data_master_writedata;                                                                      // nios2_communication:d_writedata -> nios2_communication_data_master_translator:av_writedata
	wire   [27:0] nios2_communication_data_master_address;                                                                        // nios2_communication:d_address -> nios2_communication_data_master_translator:av_address
	wire          nios2_communication_data_master_write;                                                                          // nios2_communication:d_write -> nios2_communication_data_master_translator:av_write
	wire          nios2_communication_data_master_read;                                                                           // nios2_communication:d_read -> nios2_communication_data_master_translator:av_read
	wire   [31:0] nios2_communication_data_master_readdata;                                                                       // nios2_communication_data_master_translator:av_readdata -> nios2_communication:d_readdata
	wire          nios2_communication_data_master_debugaccess;                                                                    // nios2_communication:jtag_debug_module_debugaccess_to_roms -> nios2_communication_data_master_translator:av_debugaccess
	wire    [3:0] nios2_communication_data_master_byteenable;                                                                     // nios2_communication:d_byteenable -> nios2_communication_data_master_translator:av_byteenable
	wire          nios2_car_controll_data_master_waitrequest;                                                                     // nios2_car_controll_data_master_translator:av_waitrequest -> nios2_car_controll:d_waitrequest
	wire   [31:0] nios2_car_controll_data_master_writedata;                                                                       // nios2_car_controll:d_writedata -> nios2_car_controll_data_master_translator:av_writedata
	wire   [27:0] nios2_car_controll_data_master_address;                                                                         // nios2_car_controll:d_address -> nios2_car_controll_data_master_translator:av_address
	wire          nios2_car_controll_data_master_write;                                                                           // nios2_car_controll:d_write -> nios2_car_controll_data_master_translator:av_write
	wire          nios2_car_controll_data_master_read;                                                                            // nios2_car_controll:d_read -> nios2_car_controll_data_master_translator:av_read
	wire   [31:0] nios2_car_controll_data_master_readdata;                                                                        // nios2_car_controll_data_master_translator:av_readdata -> nios2_car_controll:d_readdata
	wire          nios2_car_controll_data_master_debugaccess;                                                                     // nios2_car_controll:jtag_debug_module_debugaccess_to_roms -> nios2_car_controll_data_master_translator:av_debugaccess
	wire    [3:0] nios2_car_controll_data_master_byteenable;                                                                      // nios2_car_controll:d_byteenable -> nios2_car_controll_data_master_translator:av_byteenable
	wire          nios2_car_controll_instruction_master_waitrequest;                                                              // nios2_car_controll_instruction_master_translator:av_waitrequest -> nios2_car_controll:i_waitrequest
	wire   [18:0] nios2_car_controll_instruction_master_address;                                                                  // nios2_car_controll:i_address -> nios2_car_controll_instruction_master_translator:av_address
	wire          nios2_car_controll_instruction_master_read;                                                                     // nios2_car_controll:i_read -> nios2_car_controll_instruction_master_translator:av_read
	wire   [31:0] nios2_car_controll_instruction_master_readdata;                                                                 // nios2_car_controll_instruction_master_translator:av_readdata -> nios2_car_controll:i_readdata
	wire          nios2_car_controll_instruction_master_readdatavalid;                                                            // nios2_car_controll_instruction_master_translator:av_readdatavalid -> nios2_car_controll:i_readdatavalid
	wire          sgdma_rx_m_write_waitrequest;                                                                                   // sgdma_rx_m_write_translator:av_waitrequest -> sgdma_rx:m_write_waitrequest
	wire   [31:0] sgdma_rx_m_write_writedata;                                                                                     // sgdma_rx:m_write_writedata -> sgdma_rx_m_write_translator:av_writedata
	wire   [31:0] sgdma_rx_m_write_address;                                                                                       // sgdma_rx:m_write_address -> sgdma_rx_m_write_translator:av_address
	wire          sgdma_rx_m_write_write;                                                                                         // sgdma_rx:m_write_write -> sgdma_rx_m_write_translator:av_write
	wire    [3:0] sgdma_rx_m_write_byteenable;                                                                                    // sgdma_rx:m_write_byteenable -> sgdma_rx_m_write_translator:av_byteenable
	wire          sgdma_tx_m_read_waitrequest;                                                                                    // sgdma_tx_m_read_translator:av_waitrequest -> sgdma_tx:m_read_waitrequest
	wire   [31:0] sgdma_tx_m_read_address;                                                                                        // sgdma_tx:m_read_address -> sgdma_tx_m_read_translator:av_address
	wire          sgdma_tx_m_read_read;                                                                                           // sgdma_tx:m_read_read -> sgdma_tx_m_read_translator:av_read
	wire   [31:0] sgdma_tx_m_read_readdata;                                                                                       // sgdma_tx_m_read_translator:av_readdata -> sgdma_tx:m_read_readdata
	wire          sgdma_tx_m_read_readdatavalid;                                                                                  // sgdma_tx_m_read_translator:av_readdatavalid -> sgdma_tx:m_read_readdatavalid
	wire          sgdma_rx_descriptor_read_waitrequest;                                                                           // sgdma_rx_descriptor_read_translator:av_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	wire   [31:0] sgdma_rx_descriptor_read_address;                                                                               // sgdma_rx:descriptor_read_address -> sgdma_rx_descriptor_read_translator:av_address
	wire          sgdma_rx_descriptor_read_read;                                                                                  // sgdma_rx:descriptor_read_read -> sgdma_rx_descriptor_read_translator:av_read
	wire   [31:0] sgdma_rx_descriptor_read_readdata;                                                                              // sgdma_rx_descriptor_read_translator:av_readdata -> sgdma_rx:descriptor_read_readdata
	wire          sgdma_rx_descriptor_read_readdatavalid;                                                                         // sgdma_rx_descriptor_read_translator:av_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	wire          sgdma_rx_descriptor_write_waitrequest;                                                                          // sgdma_rx_descriptor_write_translator:av_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	wire   [31:0] sgdma_rx_descriptor_write_writedata;                                                                            // sgdma_rx:descriptor_write_writedata -> sgdma_rx_descriptor_write_translator:av_writedata
	wire   [31:0] sgdma_rx_descriptor_write_address;                                                                              // sgdma_rx:descriptor_write_address -> sgdma_rx_descriptor_write_translator:av_address
	wire          sgdma_rx_descriptor_write_write;                                                                                // sgdma_rx:descriptor_write_write -> sgdma_rx_descriptor_write_translator:av_write
	wire          sgdma_tx_descriptor_read_waitrequest;                                                                           // sgdma_tx_descriptor_read_translator:av_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	wire   [31:0] sgdma_tx_descriptor_read_address;                                                                               // sgdma_tx:descriptor_read_address -> sgdma_tx_descriptor_read_translator:av_address
	wire          sgdma_tx_descriptor_read_read;                                                                                  // sgdma_tx:descriptor_read_read -> sgdma_tx_descriptor_read_translator:av_read
	wire   [31:0] sgdma_tx_descriptor_read_readdata;                                                                              // sgdma_tx_descriptor_read_translator:av_readdata -> sgdma_tx:descriptor_read_readdata
	wire          sgdma_tx_descriptor_read_readdatavalid;                                                                         // sgdma_tx_descriptor_read_translator:av_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	wire          sgdma_tx_descriptor_write_waitrequest;                                                                          // sgdma_tx_descriptor_write_translator:av_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	wire   [31:0] sgdma_tx_descriptor_write_writedata;                                                                            // sgdma_tx:descriptor_write_writedata -> sgdma_tx_descriptor_write_translator:av_writedata
	wire   [31:0] sgdma_tx_descriptor_write_address;                                                                              // sgdma_tx:descriptor_write_address -> sgdma_tx_descriptor_write_translator:av_address
	wire          sgdma_tx_descriptor_write_write;                                                                                // sgdma_tx:descriptor_write_write -> sgdma_tx_descriptor_write_translator:av_write
	wire   [31:0] nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                 // nios2_communication_jtag_debug_module_translator:av_writedata -> nios2_communication:jtag_debug_module_writedata
	wire    [8:0] nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_address;                                   // nios2_communication_jtag_debug_module_translator:av_address -> nios2_communication:jtag_debug_module_address
	wire          nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                // nios2_communication_jtag_debug_module_translator:av_chipselect -> nios2_communication:jtag_debug_module_select
	wire          nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_write;                                     // nios2_communication_jtag_debug_module_translator:av_write -> nios2_communication:jtag_debug_module_write
	wire   [31:0] nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                  // nios2_communication:jtag_debug_module_readdata -> nios2_communication_jtag_debug_module_translator:av_readdata
	wire          nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                             // nios2_communication_jtag_debug_module_translator:av_begintransfer -> nios2_communication:jtag_debug_module_begintransfer
	wire          nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                               // nios2_communication_jtag_debug_module_translator:av_debugaccess -> nios2_communication:jtag_debug_module_debugaccess
	wire    [3:0] nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                // nios2_communication_jtag_debug_module_translator:av_byteenable -> nios2_communication:jtag_debug_module_byteenable
	wire   [31:0] main_memory_communication_s1_translator_avalon_anti_slave_0_writedata;                                          // main_memory_communication_s1_translator:av_writedata -> main_memory_communication:writedata
	wire   [14:0] main_memory_communication_s1_translator_avalon_anti_slave_0_address;                                            // main_memory_communication_s1_translator:av_address -> main_memory_communication:address
	wire          main_memory_communication_s1_translator_avalon_anti_slave_0_chipselect;                                         // main_memory_communication_s1_translator:av_chipselect -> main_memory_communication:chipselect
	wire          main_memory_communication_s1_translator_avalon_anti_slave_0_clken;                                              // main_memory_communication_s1_translator:av_clken -> main_memory_communication:clken
	wire          main_memory_communication_s1_translator_avalon_anti_slave_0_write;                                              // main_memory_communication_s1_translator:av_write -> main_memory_communication:write
	wire   [31:0] main_memory_communication_s1_translator_avalon_anti_slave_0_readdata;                                           // main_memory_communication:readdata -> main_memory_communication_s1_translator:av_readdata
	wire    [3:0] main_memory_communication_s1_translator_avalon_anti_slave_0_byteenable;                                         // main_memory_communication_s1_translator:av_byteenable -> main_memory_communication:byteenable
	wire          sdram_communication_s1_translator_avalon_anti_slave_0_waitrequest;                                              // sdram_communication:za_waitrequest -> sdram_communication_s1_translator:av_waitrequest
	wire   [31:0] sdram_communication_s1_translator_avalon_anti_slave_0_writedata;                                                // sdram_communication_s1_translator:av_writedata -> sdram_communication:az_data
	wire   [23:0] sdram_communication_s1_translator_avalon_anti_slave_0_address;                                                  // sdram_communication_s1_translator:av_address -> sdram_communication:az_addr
	wire          sdram_communication_s1_translator_avalon_anti_slave_0_chipselect;                                               // sdram_communication_s1_translator:av_chipselect -> sdram_communication:az_cs
	wire          sdram_communication_s1_translator_avalon_anti_slave_0_write;                                                    // sdram_communication_s1_translator:av_write -> sdram_communication:az_wr_n
	wire          sdram_communication_s1_translator_avalon_anti_slave_0_read;                                                     // sdram_communication_s1_translator:av_read -> sdram_communication:az_rd_n
	wire   [31:0] sdram_communication_s1_translator_avalon_anti_slave_0_readdata;                                                 // sdram_communication:za_data -> sdram_communication_s1_translator:av_readdata
	wire          sdram_communication_s1_translator_avalon_anti_slave_0_readdatavalid;                                            // sdram_communication:za_valid -> sdram_communication_s1_translator:av_readdatavalid
	wire    [3:0] sdram_communication_s1_translator_avalon_anti_slave_0_byteenable;                                               // sdram_communication_s1_translator:av_byteenable -> sdram_communication:az_be_n
	wire   [31:0] descriptor_memory_s1_translator_avalon_anti_slave_0_writedata;                                                  // descriptor_memory_s1_translator:av_writedata -> descriptor_memory:writedata
	wire    [9:0] descriptor_memory_s1_translator_avalon_anti_slave_0_address;                                                    // descriptor_memory_s1_translator:av_address -> descriptor_memory:address
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect;                                                 // descriptor_memory_s1_translator:av_chipselect -> descriptor_memory:chipselect
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_clken;                                                      // descriptor_memory_s1_translator:av_clken -> descriptor_memory:clken
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_write;                                                      // descriptor_memory_s1_translator:av_write -> descriptor_memory:write
	wire   [31:0] descriptor_memory_s1_translator_avalon_anti_slave_0_readdata;                                                   // descriptor_memory:readdata -> descriptor_memory_s1_translator:av_readdata
	wire    [3:0] descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable;                                                 // descriptor_memory_s1_translator:av_byteenable -> descriptor_memory:byteenable
	wire   [31:0] sgdma_tx_csr_translator_avalon_anti_slave_0_writedata;                                                          // sgdma_tx_csr_translator:av_writedata -> sgdma_tx:csr_writedata
	wire    [3:0] sgdma_tx_csr_translator_avalon_anti_slave_0_address;                                                            // sgdma_tx_csr_translator:av_address -> sgdma_tx:csr_address
	wire          sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect;                                                         // sgdma_tx_csr_translator:av_chipselect -> sgdma_tx:csr_chipselect
	wire          sgdma_tx_csr_translator_avalon_anti_slave_0_write;                                                              // sgdma_tx_csr_translator:av_write -> sgdma_tx:csr_write
	wire          sgdma_tx_csr_translator_avalon_anti_slave_0_read;                                                               // sgdma_tx_csr_translator:av_read -> sgdma_tx:csr_read
	wire   [31:0] sgdma_tx_csr_translator_avalon_anti_slave_0_readdata;                                                           // sgdma_tx:csr_readdata -> sgdma_tx_csr_translator:av_readdata
	wire   [31:0] sgdma_rx_csr_translator_avalon_anti_slave_0_writedata;                                                          // sgdma_rx_csr_translator:av_writedata -> sgdma_rx:csr_writedata
	wire    [3:0] sgdma_rx_csr_translator_avalon_anti_slave_0_address;                                                            // sgdma_rx_csr_translator:av_address -> sgdma_rx:csr_address
	wire          sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect;                                                         // sgdma_rx_csr_translator:av_chipselect -> sgdma_rx:csr_chipselect
	wire          sgdma_rx_csr_translator_avalon_anti_slave_0_write;                                                              // sgdma_rx_csr_translator:av_write -> sgdma_rx:csr_write
	wire          sgdma_rx_csr_translator_avalon_anti_slave_0_read;                                                               // sgdma_rx_csr_translator:av_read -> sgdma_rx:csr_read
	wire   [31:0] sgdma_rx_csr_translator_avalon_anti_slave_0_readdata;                                                           // sgdma_rx:csr_readdata -> sgdma_rx_csr_translator:av_readdata
	wire          tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest;                                                // tse_mac:waitrequest -> tse_mac_control_port_translator:av_waitrequest
	wire   [31:0] tse_mac_control_port_translator_avalon_anti_slave_0_writedata;                                                  // tse_mac_control_port_translator:av_writedata -> tse_mac:writedata
	wire    [7:0] tse_mac_control_port_translator_avalon_anti_slave_0_address;                                                    // tse_mac_control_port_translator:av_address -> tse_mac:address
	wire          tse_mac_control_port_translator_avalon_anti_slave_0_write;                                                      // tse_mac_control_port_translator:av_write -> tse_mac:write
	wire          tse_mac_control_port_translator_avalon_anti_slave_0_read;                                                       // tse_mac_control_port_translator:av_read -> tse_mac:read
	wire   [31:0] tse_mac_control_port_translator_avalon_anti_slave_0_readdata;                                                   // tse_mac:readdata -> tse_mac_control_port_translator:av_readdata
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_communication:av_waitrequest -> jtag_uart_communication_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_communication_avalon_jtag_slave_translator:av_writedata -> jtag_uart_communication:av_writedata
	wire    [0:0] jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_communication_avalon_jtag_slave_translator:av_address -> jtag_uart_communication:av_address
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_communication_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_communication:av_chipselect
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_communication_avalon_jtag_slave_translator:av_write -> jtag_uart_communication:av_write_n
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_communication_avalon_jtag_slave_translator:av_read -> jtag_uart_communication:av_read_n
	wire   [31:0] jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_communication:av_readdata -> jtag_uart_communication_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] shared_memory_s1_translator_avalon_anti_slave_0_writedata;                                                      // shared_memory_s1_translator:av_writedata -> shared_memory:writedata
	wire    [9:0] shared_memory_s1_translator_avalon_anti_slave_0_address;                                                        // shared_memory_s1_translator:av_address -> shared_memory:address
	wire          shared_memory_s1_translator_avalon_anti_slave_0_chipselect;                                                     // shared_memory_s1_translator:av_chipselect -> shared_memory:chipselect
	wire          shared_memory_s1_translator_avalon_anti_slave_0_clken;                                                          // shared_memory_s1_translator:av_clken -> shared_memory:clken
	wire          shared_memory_s1_translator_avalon_anti_slave_0_write;                                                          // shared_memory_s1_translator:av_write -> shared_memory:write
	wire   [31:0] shared_memory_s1_translator_avalon_anti_slave_0_readdata;                                                       // shared_memory:readdata -> shared_memory_s1_translator:av_readdata
	wire    [3:0] shared_memory_s1_translator_avalon_anti_slave_0_byteenable;                                                     // shared_memory_s1_translator:av_byteenable -> shared_memory:byteenable
	wire   [31:0] mutex_shared_memory_s1_translator_avalon_anti_slave_0_writedata;                                                // mutex_shared_memory_s1_translator:av_writedata -> mutex_shared_memory:data_from_cpu
	wire    [0:0] mutex_shared_memory_s1_translator_avalon_anti_slave_0_address;                                                  // mutex_shared_memory_s1_translator:av_address -> mutex_shared_memory:address
	wire          mutex_shared_memory_s1_translator_avalon_anti_slave_0_chipselect;                                               // mutex_shared_memory_s1_translator:av_chipselect -> mutex_shared_memory:chipselect
	wire          mutex_shared_memory_s1_translator_avalon_anti_slave_0_write;                                                    // mutex_shared_memory_s1_translator:av_write -> mutex_shared_memory:write
	wire          mutex_shared_memory_s1_translator_avalon_anti_slave_0_read;                                                     // mutex_shared_memory_s1_translator:av_read -> mutex_shared_memory:read
	wire   [31:0] mutex_shared_memory_s1_translator_avalon_anti_slave_0_readdata;                                                 // mutex_shared_memory:data_to_cpu -> mutex_shared_memory_s1_translator:av_readdata
	wire   [15:0] interval_timer_s1_translator_avalon_anti_slave_0_writedata;                                                     // interval_timer_s1_translator:av_writedata -> interval_timer:writedata
	wire    [2:0] interval_timer_s1_translator_avalon_anti_slave_0_address;                                                       // interval_timer_s1_translator:av_address -> interval_timer:address
	wire          interval_timer_s1_translator_avalon_anti_slave_0_chipselect;                                                    // interval_timer_s1_translator:av_chipselect -> interval_timer:chipselect
	wire          interval_timer_s1_translator_avalon_anti_slave_0_write;                                                         // interval_timer_s1_translator:av_write -> interval_timer:write_n
	wire   [15:0] interval_timer_s1_translator_avalon_anti_slave_0_readdata;                                                      // interval_timer:readdata -> interval_timer_s1_translator:av_readdata
	wire   [31:0] pio_communication_led_s1_translator_avalon_anti_slave_0_writedata;                                              // pio_communication_led_s1_translator:av_writedata -> pio_communication_led:writedata
	wire    [1:0] pio_communication_led_s1_translator_avalon_anti_slave_0_address;                                                // pio_communication_led_s1_translator:av_address -> pio_communication_led:address
	wire          pio_communication_led_s1_translator_avalon_anti_slave_0_chipselect;                                             // pio_communication_led_s1_translator:av_chipselect -> pio_communication_led:chipselect
	wire          pio_communication_led_s1_translator_avalon_anti_slave_0_write;                                                  // pio_communication_led_s1_translator:av_write -> pio_communication_led:write_n
	wire   [31:0] pio_communication_led_s1_translator_avalon_anti_slave_0_readdata;                                               // pio_communication_led:readdata -> pio_communication_led_s1_translator:av_readdata
	wire   [31:0] shared_memory_s2_translator_avalon_anti_slave_0_writedata;                                                      // shared_memory_s2_translator:av_writedata -> shared_memory:writedata2
	wire    [9:0] shared_memory_s2_translator_avalon_anti_slave_0_address;                                                        // shared_memory_s2_translator:av_address -> shared_memory:address2
	wire          shared_memory_s2_translator_avalon_anti_slave_0_chipselect;                                                     // shared_memory_s2_translator:av_chipselect -> shared_memory:chipselect2
	wire          shared_memory_s2_translator_avalon_anti_slave_0_clken;                                                          // shared_memory_s2_translator:av_clken -> shared_memory:clken2
	wire          shared_memory_s2_translator_avalon_anti_slave_0_write;                                                          // shared_memory_s2_translator:av_write -> shared_memory:write2
	wire   [31:0] shared_memory_s2_translator_avalon_anti_slave_0_readdata;                                                       // shared_memory:readdata2 -> shared_memory_s2_translator:av_readdata
	wire    [3:0] shared_memory_s2_translator_avalon_anti_slave_0_byteenable;                                                     // shared_memory_s2_translator:av_byteenable -> shared_memory:byteenable2
	wire   [31:0] main_memory_car_controll_s1_translator_avalon_anti_slave_0_writedata;                                           // main_memory_car_controll_s1_translator:av_writedata -> main_memory_car_controll:writedata
	wire   [14:0] main_memory_car_controll_s1_translator_avalon_anti_slave_0_address;                                             // main_memory_car_controll_s1_translator:av_address -> main_memory_car_controll:address
	wire          main_memory_car_controll_s1_translator_avalon_anti_slave_0_chipselect;                                          // main_memory_car_controll_s1_translator:av_chipselect -> main_memory_car_controll:chipselect
	wire          main_memory_car_controll_s1_translator_avalon_anti_slave_0_clken;                                               // main_memory_car_controll_s1_translator:av_clken -> main_memory_car_controll:clken
	wire          main_memory_car_controll_s1_translator_avalon_anti_slave_0_write;                                               // main_memory_car_controll_s1_translator:av_write -> main_memory_car_controll:write
	wire   [31:0] main_memory_car_controll_s1_translator_avalon_anti_slave_0_readdata;                                            // main_memory_car_controll:readdata -> main_memory_car_controll_s1_translator:av_readdata
	wire    [3:0] main_memory_car_controll_s1_translator_avalon_anti_slave_0_byteenable;                                          // main_memory_car_controll_s1_translator:av_byteenable -> main_memory_car_controll:byteenable
	wire   [31:0] nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                  // nios2_car_controll_jtag_debug_module_translator:av_writedata -> nios2_car_controll:jtag_debug_module_writedata
	wire    [8:0] nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_address;                                    // nios2_car_controll_jtag_debug_module_translator:av_address -> nios2_car_controll:jtag_debug_module_address
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                 // nios2_car_controll_jtag_debug_module_translator:av_chipselect -> nios2_car_controll:jtag_debug_module_select
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_write;                                      // nios2_car_controll_jtag_debug_module_translator:av_write -> nios2_car_controll:jtag_debug_module_write
	wire   [31:0] nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                   // nios2_car_controll:jtag_debug_module_readdata -> nios2_car_controll_jtag_debug_module_translator:av_readdata
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                              // nios2_car_controll_jtag_debug_module_translator:av_begintransfer -> nios2_car_controll:jtag_debug_module_begintransfer
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                // nios2_car_controll_jtag_debug_module_translator:av_debugaccess -> nios2_car_controll:jtag_debug_module_debugaccess
	wire    [3:0] nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                 // nios2_car_controll_jtag_debug_module_translator:av_byteenable -> nios2_car_controll:jtag_debug_module_byteenable
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                              // jtag_uart_carControl:av_waitrequest -> jtag_uart_carControl_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                // jtag_uart_carControl_avalon_jtag_slave_translator:av_writedata -> jtag_uart_carControl:av_writedata
	wire    [0:0] jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                  // jtag_uart_carControl_avalon_jtag_slave_translator:av_address -> jtag_uart_carControl:av_address
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                               // jtag_uart_carControl_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_carControl:av_chipselect
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                    // jtag_uart_carControl_avalon_jtag_slave_translator:av_write -> jtag_uart_carControl:av_write_n
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                     // jtag_uart_carControl_avalon_jtag_slave_translator:av_read -> jtag_uart_carControl:av_read_n
	wire   [31:0] jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                 // jtag_uart_carControl:av_readdata -> jtag_uart_carControl_avalon_jtag_slave_translator:av_readdata
	wire          nios2_communication_instruction_master_translator_avalon_universal_master_0_waitrequest;                        // nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_communication_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_communication_instruction_master_translator_avalon_universal_master_0_burstcount;                         // nios2_communication_instruction_master_translator:uav_burstcount -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_communication_instruction_master_translator_avalon_universal_master_0_writedata;                          // nios2_communication_instruction_master_translator:uav_writedata -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_communication_instruction_master_translator_avalon_universal_master_0_address;                            // nios2_communication_instruction_master_translator:uav_address -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_communication_instruction_master_translator_avalon_universal_master_0_lock;                               // nios2_communication_instruction_master_translator:uav_lock -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_communication_instruction_master_translator_avalon_universal_master_0_write;                              // nios2_communication_instruction_master_translator:uav_write -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_communication_instruction_master_translator_avalon_universal_master_0_read;                               // nios2_communication_instruction_master_translator:uav_read -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_communication_instruction_master_translator_avalon_universal_master_0_readdata;                           // nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_communication_instruction_master_translator:uav_readdata
	wire          nios2_communication_instruction_master_translator_avalon_universal_master_0_debugaccess;                        // nios2_communication_instruction_master_translator:uav_debugaccess -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_communication_instruction_master_translator_avalon_universal_master_0_byteenable;                         // nios2_communication_instruction_master_translator:uav_byteenable -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_communication_instruction_master_translator_avalon_universal_master_0_readdatavalid;                      // nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_communication_instruction_master_translator:uav_readdatavalid
	wire          nios2_communication_data_master_translator_avalon_universal_master_0_waitrequest;                               // nios2_communication_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_communication_data_master_translator:uav_waitrequest
	wire    [2:0] nios2_communication_data_master_translator_avalon_universal_master_0_burstcount;                                // nios2_communication_data_master_translator:uav_burstcount -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_communication_data_master_translator_avalon_universal_master_0_writedata;                                 // nios2_communication_data_master_translator:uav_writedata -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_communication_data_master_translator_avalon_universal_master_0_address;                                   // nios2_communication_data_master_translator:uav_address -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_communication_data_master_translator_avalon_universal_master_0_lock;                                      // nios2_communication_data_master_translator:uav_lock -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_communication_data_master_translator_avalon_universal_master_0_write;                                     // nios2_communication_data_master_translator:uav_write -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_communication_data_master_translator_avalon_universal_master_0_read;                                      // nios2_communication_data_master_translator:uav_read -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_communication_data_master_translator_avalon_universal_master_0_readdata;                                  // nios2_communication_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_communication_data_master_translator:uav_readdata
	wire          nios2_communication_data_master_translator_avalon_universal_master_0_debugaccess;                               // nios2_communication_data_master_translator:uav_debugaccess -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_communication_data_master_translator_avalon_universal_master_0_byteenable;                                // nios2_communication_data_master_translator:uav_byteenable -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_communication_data_master_translator_avalon_universal_master_0_readdatavalid;                             // nios2_communication_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_communication_data_master_translator:uav_readdatavalid
	wire          nios2_car_controll_data_master_translator_avalon_universal_master_0_waitrequest;                                // nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_car_controll_data_master_translator:uav_waitrequest
	wire    [2:0] nios2_car_controll_data_master_translator_avalon_universal_master_0_burstcount;                                 // nios2_car_controll_data_master_translator:uav_burstcount -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_car_controll_data_master_translator_avalon_universal_master_0_writedata;                                  // nios2_car_controll_data_master_translator:uav_writedata -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_car_controll_data_master_translator_avalon_universal_master_0_address;                                    // nios2_car_controll_data_master_translator:uav_address -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_car_controll_data_master_translator_avalon_universal_master_0_lock;                                       // nios2_car_controll_data_master_translator:uav_lock -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_car_controll_data_master_translator_avalon_universal_master_0_write;                                      // nios2_car_controll_data_master_translator:uav_write -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_car_controll_data_master_translator_avalon_universal_master_0_read;                                       // nios2_car_controll_data_master_translator:uav_read -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_car_controll_data_master_translator_avalon_universal_master_0_readdata;                                   // nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_car_controll_data_master_translator:uav_readdata
	wire          nios2_car_controll_data_master_translator_avalon_universal_master_0_debugaccess;                                // nios2_car_controll_data_master_translator:uav_debugaccess -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_car_controll_data_master_translator_avalon_universal_master_0_byteenable;                                 // nios2_car_controll_data_master_translator:uav_byteenable -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_car_controll_data_master_translator_avalon_universal_master_0_readdatavalid;                              // nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_car_controll_data_master_translator:uav_readdatavalid
	wire          nios2_car_controll_instruction_master_translator_avalon_universal_master_0_waitrequest;                         // nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_car_controll_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_car_controll_instruction_master_translator_avalon_universal_master_0_burstcount;                          // nios2_car_controll_instruction_master_translator:uav_burstcount -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_car_controll_instruction_master_translator_avalon_universal_master_0_writedata;                           // nios2_car_controll_instruction_master_translator:uav_writedata -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_car_controll_instruction_master_translator_avalon_universal_master_0_address;                             // nios2_car_controll_instruction_master_translator:uav_address -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_car_controll_instruction_master_translator_avalon_universal_master_0_lock;                                // nios2_car_controll_instruction_master_translator:uav_lock -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_car_controll_instruction_master_translator_avalon_universal_master_0_write;                               // nios2_car_controll_instruction_master_translator:uav_write -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_car_controll_instruction_master_translator_avalon_universal_master_0_read;                                // nios2_car_controll_instruction_master_translator:uav_read -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_car_controll_instruction_master_translator_avalon_universal_master_0_readdata;                            // nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_car_controll_instruction_master_translator:uav_readdata
	wire          nios2_car_controll_instruction_master_translator_avalon_universal_master_0_debugaccess;                         // nios2_car_controll_instruction_master_translator:uav_debugaccess -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_car_controll_instruction_master_translator_avalon_universal_master_0_byteenable;                          // nios2_car_controll_instruction_master_translator:uav_byteenable -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_car_controll_instruction_master_translator_avalon_universal_master_0_readdatavalid;                       // nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_car_controll_instruction_master_translator:uav_readdatavalid
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest;                                      // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_descriptor_read_translator:uav_waitrequest
	wire    [2:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount;                                       // sgdma_rx_descriptor_read_translator:uav_burstcount -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata;                                        // sgdma_rx_descriptor_read_translator:uav_writedata -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address;                                          // sgdma_rx_descriptor_read_translator:uav_address -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock;                                             // sgdma_rx_descriptor_read_translator:uav_lock -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write;                                            // sgdma_rx_descriptor_read_translator:uav_write -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read;                                             // sgdma_rx_descriptor_read_translator:uav_read -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata;                                         // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_descriptor_read_translator:uav_readdata
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess;                                      // sgdma_rx_descriptor_read_translator:uav_debugaccess -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable;                                       // sgdma_rx_descriptor_read_translator:uav_byteenable -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid;                                    // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_descriptor_read_translator:uav_readdatavalid
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest;                                     // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_descriptor_write_translator:uav_waitrequest
	wire    [2:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount;                                      // sgdma_rx_descriptor_write_translator:uav_burstcount -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata;                                       // sgdma_rx_descriptor_write_translator:uav_writedata -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address;                                         // sgdma_rx_descriptor_write_translator:uav_address -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock;                                            // sgdma_rx_descriptor_write_translator:uav_lock -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write;                                           // sgdma_rx_descriptor_write_translator:uav_write -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read;                                            // sgdma_rx_descriptor_write_translator:uav_read -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata;                                        // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_descriptor_write_translator:uav_readdata
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess;                                     // sgdma_rx_descriptor_write_translator:uav_debugaccess -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable;                                      // sgdma_rx_descriptor_write_translator:uav_byteenable -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid;                                   // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_descriptor_write_translator:uav_readdatavalid
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest;                                      // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_descriptor_read_translator:uav_waitrequest
	wire    [2:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount;                                       // sgdma_tx_descriptor_read_translator:uav_burstcount -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata;                                        // sgdma_tx_descriptor_read_translator:uav_writedata -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address;                                          // sgdma_tx_descriptor_read_translator:uav_address -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock;                                             // sgdma_tx_descriptor_read_translator:uav_lock -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write;                                            // sgdma_tx_descriptor_read_translator:uav_write -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read;                                             // sgdma_tx_descriptor_read_translator:uav_read -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata;                                         // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_descriptor_read_translator:uav_readdata
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess;                                      // sgdma_tx_descriptor_read_translator:uav_debugaccess -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable;                                       // sgdma_tx_descriptor_read_translator:uav_byteenable -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid;                                    // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_descriptor_read_translator:uav_readdatavalid
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest;                                     // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_descriptor_write_translator:uav_waitrequest
	wire    [2:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount;                                      // sgdma_tx_descriptor_write_translator:uav_burstcount -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata;                                       // sgdma_tx_descriptor_write_translator:uav_writedata -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address;                                         // sgdma_tx_descriptor_write_translator:uav_address -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock;                                            // sgdma_tx_descriptor_write_translator:uav_lock -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write;                                           // sgdma_tx_descriptor_write_translator:uav_write -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read;                                            // sgdma_tx_descriptor_write_translator:uav_read -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata;                                        // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_descriptor_write_translator:uav_readdata
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess;                                     // sgdma_tx_descriptor_write_translator:uav_debugaccess -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable;                                      // sgdma_tx_descriptor_write_translator:uav_byteenable -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid;                                   // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_descriptor_write_translator:uav_readdatavalid
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest;                                              // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_m_write_translator:uav_waitrequest
	wire    [2:0] sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount;                                               // sgdma_rx_m_write_translator:uav_burstcount -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_rx_m_write_translator_avalon_universal_master_0_writedata;                                                // sgdma_rx_m_write_translator:uav_writedata -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_rx_m_write_translator_avalon_universal_master_0_address;                                                  // sgdma_rx_m_write_translator:uav_address -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_lock;                                                     // sgdma_rx_m_write_translator:uav_lock -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_write;                                                    // sgdma_rx_m_write_translator:uav_write -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_read;                                                     // sgdma_rx_m_write_translator:uav_read -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_rx_m_write_translator_avalon_universal_master_0_readdata;                                                 // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_m_write_translator:uav_readdata
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess;                                              // sgdma_rx_m_write_translator:uav_debugaccess -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable;                                               // sgdma_rx_m_write_translator:uav_byteenable -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid;                                            // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_m_write_translator:uav_readdatavalid
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest;                                               // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_m_read_translator:uav_waitrequest
	wire    [2:0] sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount;                                                // sgdma_tx_m_read_translator:uav_burstcount -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_tx_m_read_translator_avalon_universal_master_0_writedata;                                                 // sgdma_tx_m_read_translator:uav_writedata -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_tx_m_read_translator_avalon_universal_master_0_address;                                                   // sgdma_tx_m_read_translator:uav_address -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_lock;                                                      // sgdma_tx_m_read_translator:uav_lock -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_write;                                                     // sgdma_tx_m_read_translator:uav_write -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_read;                                                      // sgdma_tx_m_read_translator:uav_read -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_tx_m_read_translator_avalon_universal_master_0_readdata;                                                  // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_m_read_translator:uav_readdata
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess;                                               // sgdma_tx_m_read_translator:uav_debugaccess -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable;                                                // sgdma_tx_m_read_translator:uav_byteenable -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid;                                             // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_m_read_translator:uav_readdatavalid
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // nios2_communication_jtag_debug_module_translator:uav_waitrequest -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_communication_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                   // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_communication_jtag_debug_module_translator:uav_writedata
	wire   [31:0] nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                     // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_communication_jtag_debug_module_translator:uav_address
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                       // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_communication_jtag_debug_module_translator:uav_write
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                        // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_communication_jtag_debug_module_translator:uav_lock
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                        // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_communication_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                    // nios2_communication_jtag_debug_module_translator:uav_readdata -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // nios2_communication_jtag_debug_module_translator:uav_readdatavalid -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_communication_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_communication_jtag_debug_module_translator:uav_byteenable
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                 // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // main_memory_communication_s1_translator:uav_waitrequest -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> main_memory_communication_s1_translator:uav_burstcount
	wire   [31:0] main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> main_memory_communication_s1_translator:uav_writedata
	wire   [31:0] main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:m0_address -> main_memory_communication_s1_translator:uav_address
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:m0_write -> main_memory_communication_s1_translator:uav_write
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:m0_lock -> main_memory_communication_s1_translator:uav_lock
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:m0_read -> main_memory_communication_s1_translator:uav_read
	wire   [31:0] main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // main_memory_communication_s1_translator:uav_readdata -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // main_memory_communication_s1_translator:uav_readdatavalid -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> main_memory_communication_s1_translator:uav_debugaccess
	wire    [3:0] main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> main_memory_communication_s1_translator:uav_byteenable
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // sdram_communication_s1_translator:uav_waitrequest -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // sdram_communication_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_communication_s1_translator:uav_burstcount
	wire   [31:0] sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // sdram_communication_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_communication_s1_translator:uav_writedata
	wire   [31:0] sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // sdram_communication_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_communication_s1_translator:uav_address
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // sdram_communication_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_communication_s1_translator:uav_write
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // sdram_communication_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_communication_s1_translator:uav_lock
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // sdram_communication_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_communication_s1_translator:uav_read
	wire   [31:0] sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // sdram_communication_s1_translator:uav_readdata -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // sdram_communication_s1_translator:uav_readdatavalid -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // sdram_communication_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_communication_s1_translator:uav_debugaccess
	wire    [3:0] sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // sdram_communication_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_communication_s1_translator:uav_byteenable
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // sdram_communication_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // sdram_communication_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // sdram_communication_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // sdram_communication_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // sdram_communication_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // sdram_communication_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sdram_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // sdram_communication_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // sdram_communication_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // descriptor_memory_s1_translator:uav_waitrequest -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> descriptor_memory_s1_translator:uav_burstcount
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> descriptor_memory_s1_translator:uav_writedata
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> descriptor_memory_s1_translator:uav_address
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> descriptor_memory_s1_translator:uav_write
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> descriptor_memory_s1_translator:uav_lock
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> descriptor_memory_s1_translator:uav_read
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // descriptor_memory_s1_translator:uav_readdata -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // descriptor_memory_s1_translator:uav_readdatavalid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> descriptor_memory_s1_translator:uav_debugaccess
	wire    [3:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> descriptor_memory_s1_translator:uav_byteenable
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                          // sgdma_tx_csr_translator:uav_waitrequest -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                                           // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_tx_csr_translator:uav_burstcount
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                            // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_tx_csr_translator:uav_writedata
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address;                                              // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_tx_csr_translator:uav_address
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write;                                                // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_tx_csr_translator:uav_write
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_tx_csr_translator:uav_lock
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read;                                                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_tx_csr_translator:uav_read
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                             // sgdma_tx_csr_translator:uav_readdata -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                        // sgdma_tx_csr_translator:uav_readdatavalid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                          // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_tx_csr_translator:uav_debugaccess
	wire    [3:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                                           // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_tx_csr_translator:uav_byteenable
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                   // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                                         // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                                          // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                                         // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                      // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                              // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                       // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                      // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                    // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                     // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                    // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                          // sgdma_rx_csr_translator:uav_waitrequest -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                                           // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_rx_csr_translator:uav_burstcount
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                            // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_rx_csr_translator:uav_writedata
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address;                                              // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_rx_csr_translator:uav_address
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write;                                                // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_rx_csr_translator:uav_write
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_rx_csr_translator:uav_lock
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read;                                                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_rx_csr_translator:uav_read
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                             // sgdma_rx_csr_translator:uav_readdata -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                        // sgdma_rx_csr_translator:uav_readdatavalid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                          // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_rx_csr_translator:uav_debugaccess
	wire    [3:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                                           // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_rx_csr_translator:uav_byteenable
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                   // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                                         // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                                          // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                                         // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                      // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                              // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                       // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                      // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                    // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                     // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                    // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // tse_mac_control_port_translator:uav_waitrequest -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> tse_mac_control_port_translator:uav_burstcount
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> tse_mac_control_port_translator:uav_writedata
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address;                                      // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_address -> tse_mac_control_port_translator:uav_address
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write;                                        // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_write -> tse_mac_control_port_translator:uav_write
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                                         // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> tse_mac_control_port_translator:uav_lock
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read;                                         // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_read -> tse_mac_control_port_translator:uav_read
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // tse_mac_control_port_translator:uav_readdata -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // tse_mac_control_port_translator:uav_readdatavalid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> tse_mac_control_port_translator:uav_debugaccess
	wire    [3:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> tse_mac_control_port_translator:uav_byteenable
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_communication_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_communication_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_communication_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_communication_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_communication_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_communication_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_communication_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_communication_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_communication_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_communication_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_communication_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // shared_memory_s1_translator:uav_waitrequest -> shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> shared_memory_s1_translator:uav_burstcount
	wire   [31:0] shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> shared_memory_s1_translator:uav_writedata
	wire   [31:0] shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> shared_memory_s1_translator:uav_address
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> shared_memory_s1_translator:uav_write
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> shared_memory_s1_translator:uav_lock
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> shared_memory_s1_translator:uav_read
	wire   [31:0] shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // shared_memory_s1_translator:uav_readdata -> shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // shared_memory_s1_translator:uav_readdatavalid -> shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> shared_memory_s1_translator:uav_debugaccess
	wire    [3:0] shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> shared_memory_s1_translator:uav_byteenable
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // shared_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> shared_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // shared_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> shared_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // shared_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> shared_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // mutex_shared_memory_s1_translator:uav_waitrequest -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> mutex_shared_memory_s1_translator:uav_burstcount
	wire   [31:0] mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> mutex_shared_memory_s1_translator:uav_writedata
	wire   [31:0] mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> mutex_shared_memory_s1_translator:uav_address
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> mutex_shared_memory_s1_translator:uav_write
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> mutex_shared_memory_s1_translator:uav_lock
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> mutex_shared_memory_s1_translator:uav_read
	wire   [31:0] mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // mutex_shared_memory_s1_translator:uav_readdata -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // mutex_shared_memory_s1_translator:uav_readdatavalid -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mutex_shared_memory_s1_translator:uav_debugaccess
	wire    [3:0] mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> mutex_shared_memory_s1_translator:uav_byteenable
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // interval_timer_s1_translator:uav_waitrequest -> interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> interval_timer_s1_translator:uav_burstcount
	wire   [31:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> interval_timer_s1_translator:uav_writedata
	wire   [31:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> interval_timer_s1_translator:uav_address
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> interval_timer_s1_translator:uav_write
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> interval_timer_s1_translator:uav_lock
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> interval_timer_s1_translator:uav_read
	wire   [31:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // interval_timer_s1_translator:uav_readdata -> interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // interval_timer_s1_translator:uav_readdatavalid -> interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> interval_timer_s1_translator:uav_debugaccess
	wire    [3:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> interval_timer_s1_translator:uav_byteenable
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // pio_communication_led_s1_translator:uav_waitrequest -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_communication_led_s1_translator:uav_burstcount
	wire   [31:0] pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_communication_led_s1_translator:uav_writedata
	wire   [31:0] pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_communication_led_s1_translator:uav_address
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_communication_led_s1_translator:uav_write
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_communication_led_s1_translator:uav_lock
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_communication_led_s1_translator:uav_read
	wire   [31:0] pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // pio_communication_led_s1_translator:uav_readdata -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // pio_communication_led_s1_translator:uav_readdatavalid -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_communication_led_s1_translator:uav_debugaccess
	wire    [3:0] pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_communication_led_s1_translator:uav_byteenable
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // shared_memory_s2_translator:uav_waitrequest -> shared_memory_s2_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // shared_memory_s2_translator_avalon_universal_slave_0_agent:m0_burstcount -> shared_memory_s2_translator:uav_burstcount
	wire   [31:0] shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // shared_memory_s2_translator_avalon_universal_slave_0_agent:m0_writedata -> shared_memory_s2_translator:uav_writedata
	wire   [31:0] shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_address;                                          // shared_memory_s2_translator_avalon_universal_slave_0_agent:m0_address -> shared_memory_s2_translator:uav_address
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_write;                                            // shared_memory_s2_translator_avalon_universal_slave_0_agent:m0_write -> shared_memory_s2_translator:uav_write
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_lock;                                             // shared_memory_s2_translator_avalon_universal_slave_0_agent:m0_lock -> shared_memory_s2_translator:uav_lock
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_read;                                             // shared_memory_s2_translator_avalon_universal_slave_0_agent:m0_read -> shared_memory_s2_translator:uav_read
	wire   [31:0] shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // shared_memory_s2_translator:uav_readdata -> shared_memory_s2_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // shared_memory_s2_translator:uav_readdatavalid -> shared_memory_s2_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // shared_memory_s2_translator_avalon_universal_slave_0_agent:m0_debugaccess -> shared_memory_s2_translator:uav_debugaccess
	wire    [3:0] shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // shared_memory_s2_translator_avalon_universal_slave_0_agent:m0_byteenable -> shared_memory_s2_translator:uav_byteenable
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // shared_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // shared_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_valid -> shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // shared_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // shared_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_data -> shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> shared_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> shared_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> shared_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> shared_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> shared_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // shared_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_ready -> shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // shared_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> shared_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] shared_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // shared_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> shared_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // shared_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> shared_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // main_memory_car_controll_s1_translator:uav_waitrequest -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> main_memory_car_controll_s1_translator:uav_burstcount
	wire   [31:0] main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> main_memory_car_controll_s1_translator:uav_writedata
	wire   [31:0] main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:m0_address -> main_memory_car_controll_s1_translator:uav_address
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:m0_write -> main_memory_car_controll_s1_translator:uav_write
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:m0_lock -> main_memory_car_controll_s1_translator:uav_lock
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:m0_read -> main_memory_car_controll_s1_translator:uav_read
	wire   [31:0] main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // main_memory_car_controll_s1_translator:uav_readdata -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // main_memory_car_controll_s1_translator:uav_readdatavalid -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> main_memory_car_controll_s1_translator:uav_debugaccess
	wire    [3:0] main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> main_memory_car_controll_s1_translator:uav_byteenable
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // nios2_car_controll_jtag_debug_module_translator:uav_waitrequest -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_car_controll_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                    // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_car_controll_jtag_debug_module_translator:uav_writedata
	wire   [31:0] nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                      // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_car_controll_jtag_debug_module_translator:uav_address
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                        // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_car_controll_jtag_debug_module_translator:uav_write
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                         // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_car_controll_jtag_debug_module_translator:uav_lock
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                         // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_car_controll_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                     // nios2_car_controll_jtag_debug_module_translator:uav_readdata -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // nios2_car_controll_jtag_debug_module_translator:uav_readdatavalid -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_car_controll_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_car_controll_jtag_debug_module_translator:uav_byteenable
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                  // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // jtag_uart_carControl_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_carControl_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_carControl_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_carControl_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_carControl_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_carControl_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_carControl_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // jtag_uart_carControl_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // jtag_uart_carControl_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_carControl_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_carControl_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;               // nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                     // nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;             // nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [106:0] nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                      // nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router:sink_ready -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // nios2_communication_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_valid;                            // nios2_communication_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // nios2_communication_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [106:0] nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_data;                             // nios2_communication_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_001:sink_ready -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_valid;                             // nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [106:0] nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_data;                              // nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_002:sink_ready -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                // nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                      // nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;              // nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [106:0] nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                       // nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                      // addr_router_003:sink_ready -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                             // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;                                   // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                           // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [106:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;                                    // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;                                   // addr_router_004:sink_ready -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                            // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;                                  // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;                          // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire  [106:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;                                   // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;                                  // addr_router_005:sink_ready -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                             // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_006:sink_endofpacket
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;                                   // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_006:sink_valid
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                           // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_006:sink_startofpacket
	wire  [106:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;                                    // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_006:sink_data
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;                                   // addr_router_006:sink_ready -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                            // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_007:sink_endofpacket
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;                                  // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_007:sink_valid
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;                          // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_007:sink_startofpacket
	wire  [106:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;                                   // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_007:sink_data
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;                                  // addr_router_007:sink_ready -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                                     // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_008:sink_endofpacket
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid;                                           // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_008:sink_valid
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket;                                   // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_008:sink_startofpacket
	wire  [106:0] sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data;                                            // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_008:sink_data
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready;                                           // addr_router_008:sink_ready -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                                      // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_009:sink_endofpacket
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid;                                            // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_009:sink_valid
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                                    // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_009:sink_startofpacket
	wire  [106:0] sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data;                                             // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_009:sink_data
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready;                                            // addr_router_009:sink_ready -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                       // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [106:0] nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                        // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router:sink_ready -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [106:0] main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_001:sink_ready -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // sdram_communication_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // sdram_communication_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // sdram_communication_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [106:0] sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // sdram_communication_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_002:sink_ready -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [106:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_003:sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                          // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                                // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                        // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [106:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data;                                                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                                // id_router_004:sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                          // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                                // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                        // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [106:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data;                                                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                                // id_router_005:sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                                        // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [106:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data;                                         // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_006:sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [106:0] jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_007:sink_ready -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // shared_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // shared_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // shared_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [106:0] shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // shared_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_008:sink_ready -> shared_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [106:0] mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_009:sink_ready -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [106:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_010:sink_ready -> interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [106:0] pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_011:sink_ready -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // shared_memory_s2_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_valid;                                            // shared_memory_s2_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // shared_memory_s2_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [106:0] shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_data;                                             // shared_memory_s2_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_012:sink_ready -> shared_memory_s2_translator_avalon_universal_slave_0_agent:rp_ready
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [106:0] main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_013:sink_ready -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                        // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [106:0] nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                         // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_014:sink_ready -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [106:0] jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_015:sink_ready -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                                    // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                          // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                                  // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [106:0] addr_router_src_data;                                                                                           // addr_router:src_data -> limiter:cmd_sink_data
	wire   [15:0] addr_router_src_channel;                                                                                        // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                          // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                                    // limiter:rsp_src_endofpacket -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                          // limiter:rsp_src_valid -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                                  // limiter:rsp_src_startofpacket -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_rsp_src_data;                                                                                           // limiter:rsp_src_data -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] limiter_rsp_src_channel;                                                                                        // limiter:rsp_src_channel -> nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                          // nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_003_src_endofpacket;                                                                                // addr_router_003:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_003_src_valid;                                                                                      // addr_router_003:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_003_src_startofpacket;                                                                              // addr_router_003:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [106:0] addr_router_003_src_data;                                                                                       // addr_router_003:src_data -> limiter_001:cmd_sink_data
	wire   [15:0] addr_router_003_src_channel;                                                                                    // addr_router_003:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_003_src_ready;                                                                                      // limiter_001:cmd_sink_ready -> addr_router_003:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                                // limiter_001:rsp_src_endofpacket -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                                      // limiter_001:rsp_src_valid -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                              // limiter_001:rsp_src_startofpacket -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_001_rsp_src_data;                                                                                       // limiter_001:rsp_src_data -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] limiter_001_rsp_src_channel;                                                                                    // limiter_001:rsp_src_channel -> nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                                      // nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          rst_controller_reset_out_reset;                                                                                 // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, addr_router_005:reset, addr_router_006:reset, addr_router_007:reset, addr_router_008:reset, addr_router_009:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_demux_005:reset, cmd_xbar_demux_006:reset, cmd_xbar_demux_007:reset, cmd_xbar_demux_008:reset, cmd_xbar_demux_009:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_009:reset, cmd_xbar_mux_010:reset, cmd_xbar_mux_013:reset, cmd_xbar_mux_014:reset, descriptor_memory:reset, descriptor_memory_s1_translator:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, interval_timer:reset_n, interval_timer_s1_translator:reset, interval_timer_s1_translator_avalon_universal_slave_0_agent:reset, interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, irq_mapper:reset, irq_mapper_001:reset, jtag_uart_carControl:rst_n, jtag_uart_carControl_avalon_jtag_slave_translator:reset, jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, jtag_uart_communication:rst_n, jtag_uart_communication_avalon_jtag_slave_translator:reset, jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, main_memory_car_controll:reset, main_memory_car_controll_s1_translator:reset, main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:reset, main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, main_memory_communication:reset, main_memory_communication_s1_translator:reset, main_memory_communication_s1_translator_avalon_universal_slave_0_agent:reset, main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mutex_shared_memory:reset_n, mutex_shared_memory_s1_translator:reset, mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:reset, mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_car_controll:reset_n, nios2_car_controll_data_master_translator:reset, nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:reset, nios2_car_controll_instruction_master_translator:reset, nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_car_controll_jtag_debug_module_translator:reset, nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_communication:reset_n, nios2_communication_data_master_translator:reset, nios2_communication_data_master_translator_avalon_universal_master_0_agent:reset, nios2_communication_instruction_master_translator:reset, nios2_communication_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_communication_jtag_debug_module_translator:reset, nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_communication_led:reset_n, pio_communication_led_s1_translator:reset, pio_communication_led_s1_translator_avalon_universal_slave_0_agent:reset, pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_002:reset, rsp_xbar_mux_003:reset, sgdma_rx:system_reset_n, sgdma_rx_csr_translator:reset, sgdma_rx_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_rx_descriptor_read_translator:reset, sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_rx_descriptor_write_translator:reset, sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_rx_m_write_translator:reset, sgdma_rx_m_write_translator_avalon_universal_master_0_agent:reset, sgdma_tx:system_reset_n, sgdma_tx_csr_translator:reset, sgdma_tx_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_tx_descriptor_read_translator:reset, sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_tx_descriptor_write_translator:reset, sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_tx_m_read_translator:reset, sgdma_tx_m_read_translator_avalon_universal_master_0_agent:reset, shared_memory:reset, shared_memory_s1_translator:reset, shared_memory_s1_translator_avalon_universal_slave_0_agent:reset, shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, shared_memory_s2_translator:reset, shared_memory_s2_translator_avalon_universal_slave_0_agent:reset, shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, tse_mac:reset, tse_mac_control_port_translator:reset, tse_mac_control_port_translator_avalon_universal_slave_0_agent:reset, tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          nios2_communication_jtag_debug_module_reset_reset;                                                              // nios2_communication:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire          nios2_car_controll_jtag_debug_module_reset_reset;                                                               // nios2_car_controll:jtag_debug_module_resetrequest -> rst_controller:reset_in2
	wire          rst_controller_001_reset_out_reset;                                                                             // rst_controller_001:reset_out -> [cmd_xbar_mux_002:reset, id_router_002:reset, rsp_xbar_demux_002:reset, sdram_communication:reset_n, sdram_communication_s1_translator:reset, sdram_communication_s1_translator_avalon_universal_slave_0_agent:reset, sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                                // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                      // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                              // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src0_data;                                                                                       // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [15:0] cmd_xbar_demux_src0_channel;                                                                                    // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                      // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                                // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                      // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                              // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src1_data;                                                                                       // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [15:0] cmd_xbar_demux_src1_channel;                                                                                    // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                      // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                                // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                      // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                              // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src2_data;                                                                                       // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [15:0] cmd_xbar_demux_src2_channel;                                                                                    // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                                      // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                            // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                  // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                          // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src0_data;                                                                                   // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [15:0] cmd_xbar_demux_001_src0_channel;                                                                                // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                                  // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                            // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                                  // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                          // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src1_data;                                                                                   // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [15:0] cmd_xbar_demux_001_src1_channel;                                                                                // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                                  // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                            // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                                  // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                          // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src2_data;                                                                                   // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [15:0] cmd_xbar_demux_001_src2_channel;                                                                                // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                                  // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                            // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                                  // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                          // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src3_data;                                                                                   // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [15:0] cmd_xbar_demux_001_src3_channel;                                                                                // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                                  // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                            // cmd_xbar_demux_001:src4_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                                  // cmd_xbar_demux_001:src4_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                          // cmd_xbar_demux_001:src4_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src4_data;                                                                                   // cmd_xbar_demux_001:src4_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src4_channel;                                                                                // cmd_xbar_demux_001:src4_channel -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                            // cmd_xbar_demux_001:src5_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                                  // cmd_xbar_demux_001:src5_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                          // cmd_xbar_demux_001:src5_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src5_data;                                                                                   // cmd_xbar_demux_001:src5_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src5_channel;                                                                                // cmd_xbar_demux_001:src5_channel -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                            // cmd_xbar_demux_001:src6_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                                  // cmd_xbar_demux_001:src6_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                          // cmd_xbar_demux_001:src6_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src6_data;                                                                                   // cmd_xbar_demux_001:src6_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src6_channel;                                                                                // cmd_xbar_demux_001:src6_channel -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                            // cmd_xbar_demux_001:src7_endofpacket -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                                  // cmd_xbar_demux_001:src7_valid -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                          // cmd_xbar_demux_001:src7_startofpacket -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src7_data;                                                                                   // cmd_xbar_demux_001:src7_data -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src7_channel;                                                                                // cmd_xbar_demux_001:src7_channel -> jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                            // cmd_xbar_demux_001:src8_endofpacket -> shared_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                                  // cmd_xbar_demux_001:src8_valid -> shared_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                          // cmd_xbar_demux_001:src8_startofpacket -> shared_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src8_data;                                                                                   // cmd_xbar_demux_001:src8_data -> shared_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src8_channel;                                                                                // cmd_xbar_demux_001:src8_channel -> shared_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                            // cmd_xbar_demux_001:src9_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                                  // cmd_xbar_demux_001:src9_valid -> cmd_xbar_mux_009:sink0_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                          // cmd_xbar_demux_001:src9_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src9_data;                                                                                   // cmd_xbar_demux_001:src9_data -> cmd_xbar_mux_009:sink0_data
	wire   [15:0] cmd_xbar_demux_001_src9_channel;                                                                                // cmd_xbar_demux_001:src9_channel -> cmd_xbar_mux_009:sink0_channel
	wire          cmd_xbar_demux_001_src9_ready;                                                                                  // cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux_001:src9_ready
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                           // cmd_xbar_demux_001:src10_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                                 // cmd_xbar_demux_001:src10_valid -> cmd_xbar_mux_010:sink0_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                         // cmd_xbar_demux_001:src10_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src10_data;                                                                                  // cmd_xbar_demux_001:src10_data -> cmd_xbar_mux_010:sink0_data
	wire   [15:0] cmd_xbar_demux_001_src10_channel;                                                                               // cmd_xbar_demux_001:src10_channel -> cmd_xbar_mux_010:sink0_channel
	wire          cmd_xbar_demux_001_src10_ready;                                                                                 // cmd_xbar_mux_010:sink0_ready -> cmd_xbar_demux_001:src10_ready
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                                           // cmd_xbar_demux_001:src11_endofpacket -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                                 // cmd_xbar_demux_001:src11_valid -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                                         // cmd_xbar_demux_001:src11_startofpacket -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src11_data;                                                                                  // cmd_xbar_demux_001:src11_data -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src11_channel;                                                                               // cmd_xbar_demux_001:src11_channel -> pio_communication_led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                            // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                                  // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_009:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                          // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src0_data;                                                                                   // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_009:sink1_data
	wire   [15:0] cmd_xbar_demux_002_src0_channel;                                                                                // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_009:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                                  // cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_002_src1_endofpacket;                                                                            // cmd_xbar_demux_002:src1_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	wire          cmd_xbar_demux_002_src1_valid;                                                                                  // cmd_xbar_demux_002:src1_valid -> cmd_xbar_mux_010:sink1_valid
	wire          cmd_xbar_demux_002_src1_startofpacket;                                                                          // cmd_xbar_demux_002:src1_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src1_data;                                                                                   // cmd_xbar_demux_002:src1_data -> cmd_xbar_mux_010:sink1_data
	wire   [15:0] cmd_xbar_demux_002_src1_channel;                                                                                // cmd_xbar_demux_002:src1_channel -> cmd_xbar_mux_010:sink1_channel
	wire          cmd_xbar_demux_002_src1_ready;                                                                                  // cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_002:src1_ready
	wire          cmd_xbar_demux_002_src2_endofpacket;                                                                            // cmd_xbar_demux_002:src2_endofpacket -> shared_memory_s2_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src2_valid;                                                                                  // cmd_xbar_demux_002:src2_valid -> shared_memory_s2_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src2_startofpacket;                                                                          // cmd_xbar_demux_002:src2_startofpacket -> shared_memory_s2_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src2_data;                                                                                   // cmd_xbar_demux_002:src2_data -> shared_memory_s2_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_002_src2_channel;                                                                                // cmd_xbar_demux_002:src2_channel -> shared_memory_s2_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src3_endofpacket;                                                                            // cmd_xbar_demux_002:src3_endofpacket -> cmd_xbar_mux_013:sink0_endofpacket
	wire          cmd_xbar_demux_002_src3_valid;                                                                                  // cmd_xbar_demux_002:src3_valid -> cmd_xbar_mux_013:sink0_valid
	wire          cmd_xbar_demux_002_src3_startofpacket;                                                                          // cmd_xbar_demux_002:src3_startofpacket -> cmd_xbar_mux_013:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src3_data;                                                                                   // cmd_xbar_demux_002:src3_data -> cmd_xbar_mux_013:sink0_data
	wire   [15:0] cmd_xbar_demux_002_src3_channel;                                                                                // cmd_xbar_demux_002:src3_channel -> cmd_xbar_mux_013:sink0_channel
	wire          cmd_xbar_demux_002_src3_ready;                                                                                  // cmd_xbar_mux_013:sink0_ready -> cmd_xbar_demux_002:src3_ready
	wire          cmd_xbar_demux_002_src4_endofpacket;                                                                            // cmd_xbar_demux_002:src4_endofpacket -> cmd_xbar_mux_014:sink0_endofpacket
	wire          cmd_xbar_demux_002_src4_valid;                                                                                  // cmd_xbar_demux_002:src4_valid -> cmd_xbar_mux_014:sink0_valid
	wire          cmd_xbar_demux_002_src4_startofpacket;                                                                          // cmd_xbar_demux_002:src4_startofpacket -> cmd_xbar_mux_014:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src4_data;                                                                                   // cmd_xbar_demux_002:src4_data -> cmd_xbar_mux_014:sink0_data
	wire   [15:0] cmd_xbar_demux_002_src4_channel;                                                                                // cmd_xbar_demux_002:src4_channel -> cmd_xbar_mux_014:sink0_channel
	wire          cmd_xbar_demux_002_src4_ready;                                                                                  // cmd_xbar_mux_014:sink0_ready -> cmd_xbar_demux_002:src4_ready
	wire          cmd_xbar_demux_002_src5_endofpacket;                                                                            // cmd_xbar_demux_002:src5_endofpacket -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_002_src5_valid;                                                                                  // cmd_xbar_demux_002:src5_valid -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_002_src5_startofpacket;                                                                          // cmd_xbar_demux_002:src5_startofpacket -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src5_data;                                                                                   // cmd_xbar_demux_002:src5_data -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_002_src5_channel;                                                                                // cmd_xbar_demux_002:src5_channel -> jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                            // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_013:sink1_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                                  // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_013:sink1_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                                          // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_013:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src0_data;                                                                                   // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_013:sink1_data
	wire   [15:0] cmd_xbar_demux_003_src0_channel;                                                                                // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_013:sink1_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                                  // cmd_xbar_mux_013:sink1_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_003_src1_endofpacket;                                                                            // cmd_xbar_demux_003:src1_endofpacket -> cmd_xbar_mux_014:sink1_endofpacket
	wire          cmd_xbar_demux_003_src1_valid;                                                                                  // cmd_xbar_demux_003:src1_valid -> cmd_xbar_mux_014:sink1_valid
	wire          cmd_xbar_demux_003_src1_startofpacket;                                                                          // cmd_xbar_demux_003:src1_startofpacket -> cmd_xbar_mux_014:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src1_data;                                                                                   // cmd_xbar_demux_003:src1_data -> cmd_xbar_mux_014:sink1_data
	wire   [15:0] cmd_xbar_demux_003_src1_channel;                                                                                // cmd_xbar_demux_003:src1_channel -> cmd_xbar_mux_014:sink1_channel
	wire          cmd_xbar_demux_003_src1_ready;                                                                                  // cmd_xbar_mux_014:sink1_ready -> cmd_xbar_demux_003:src1_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                            // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                                  // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                                          // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_004_src0_data;                                                                                   // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_003:sink1_data
	wire   [15:0] cmd_xbar_demux_004_src0_channel;                                                                                // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                                  // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_004:src0_ready
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                                            // cmd_xbar_demux_005:src0_endofpacket -> cmd_xbar_mux_003:sink2_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                                  // cmd_xbar_demux_005:src0_valid -> cmd_xbar_mux_003:sink2_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                                          // cmd_xbar_demux_005:src0_startofpacket -> cmd_xbar_mux_003:sink2_startofpacket
	wire  [106:0] cmd_xbar_demux_005_src0_data;                                                                                   // cmd_xbar_demux_005:src0_data -> cmd_xbar_mux_003:sink2_data
	wire   [15:0] cmd_xbar_demux_005_src0_channel;                                                                                // cmd_xbar_demux_005:src0_channel -> cmd_xbar_mux_003:sink2_channel
	wire          cmd_xbar_demux_005_src0_ready;                                                                                  // cmd_xbar_mux_003:sink2_ready -> cmd_xbar_demux_005:src0_ready
	wire          cmd_xbar_demux_006_src0_endofpacket;                                                                            // cmd_xbar_demux_006:src0_endofpacket -> cmd_xbar_mux_003:sink3_endofpacket
	wire          cmd_xbar_demux_006_src0_valid;                                                                                  // cmd_xbar_demux_006:src0_valid -> cmd_xbar_mux_003:sink3_valid
	wire          cmd_xbar_demux_006_src0_startofpacket;                                                                          // cmd_xbar_demux_006:src0_startofpacket -> cmd_xbar_mux_003:sink3_startofpacket
	wire  [106:0] cmd_xbar_demux_006_src0_data;                                                                                   // cmd_xbar_demux_006:src0_data -> cmd_xbar_mux_003:sink3_data
	wire   [15:0] cmd_xbar_demux_006_src0_channel;                                                                                // cmd_xbar_demux_006:src0_channel -> cmd_xbar_mux_003:sink3_channel
	wire          cmd_xbar_demux_006_src0_ready;                                                                                  // cmd_xbar_mux_003:sink3_ready -> cmd_xbar_demux_006:src0_ready
	wire          cmd_xbar_demux_007_src0_endofpacket;                                                                            // cmd_xbar_demux_007:src0_endofpacket -> cmd_xbar_mux_003:sink4_endofpacket
	wire          cmd_xbar_demux_007_src0_valid;                                                                                  // cmd_xbar_demux_007:src0_valid -> cmd_xbar_mux_003:sink4_valid
	wire          cmd_xbar_demux_007_src0_startofpacket;                                                                          // cmd_xbar_demux_007:src0_startofpacket -> cmd_xbar_mux_003:sink4_startofpacket
	wire  [106:0] cmd_xbar_demux_007_src0_data;                                                                                   // cmd_xbar_demux_007:src0_data -> cmd_xbar_mux_003:sink4_data
	wire   [15:0] cmd_xbar_demux_007_src0_channel;                                                                                // cmd_xbar_demux_007:src0_channel -> cmd_xbar_mux_003:sink4_channel
	wire          cmd_xbar_demux_007_src0_ready;                                                                                  // cmd_xbar_mux_003:sink4_ready -> cmd_xbar_demux_007:src0_ready
	wire          cmd_xbar_demux_008_src0_endofpacket;                                                                            // cmd_xbar_demux_008:src0_endofpacket -> cmd_xbar_mux_001:sink2_endofpacket
	wire          cmd_xbar_demux_008_src0_valid;                                                                                  // cmd_xbar_demux_008:src0_valid -> cmd_xbar_mux_001:sink2_valid
	wire          cmd_xbar_demux_008_src0_startofpacket;                                                                          // cmd_xbar_demux_008:src0_startofpacket -> cmd_xbar_mux_001:sink2_startofpacket
	wire  [106:0] cmd_xbar_demux_008_src0_data;                                                                                   // cmd_xbar_demux_008:src0_data -> cmd_xbar_mux_001:sink2_data
	wire   [15:0] cmd_xbar_demux_008_src0_channel;                                                                                // cmd_xbar_demux_008:src0_channel -> cmd_xbar_mux_001:sink2_channel
	wire          cmd_xbar_demux_008_src0_ready;                                                                                  // cmd_xbar_mux_001:sink2_ready -> cmd_xbar_demux_008:src0_ready
	wire          cmd_xbar_demux_009_src0_endofpacket;                                                                            // cmd_xbar_demux_009:src0_endofpacket -> cmd_xbar_mux_001:sink3_endofpacket
	wire          cmd_xbar_demux_009_src0_valid;                                                                                  // cmd_xbar_demux_009:src0_valid -> cmd_xbar_mux_001:sink3_valid
	wire          cmd_xbar_demux_009_src0_startofpacket;                                                                          // cmd_xbar_demux_009:src0_startofpacket -> cmd_xbar_mux_001:sink3_startofpacket
	wire  [106:0] cmd_xbar_demux_009_src0_data;                                                                                   // cmd_xbar_demux_009:src0_data -> cmd_xbar_mux_001:sink3_data
	wire   [15:0] cmd_xbar_demux_009_src0_channel;                                                                                // cmd_xbar_demux_009:src0_channel -> cmd_xbar_mux_001:sink3_channel
	wire          cmd_xbar_demux_009_src0_ready;                                                                                  // cmd_xbar_mux_001:sink3_ready -> cmd_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                                // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                      // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                              // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src0_data;                                                                                       // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [15:0] rsp_xbar_demux_src0_channel;                                                                                    // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                      // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                                // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                      // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                              // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src1_data;                                                                                       // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [15:0] rsp_xbar_demux_src1_channel;                                                                                    // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                      // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                            // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                  // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                          // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src0_data;                                                                                   // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [15:0] rsp_xbar_demux_001_src0_channel;                                                                                // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                  // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                            // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                                  // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                          // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src1_data;                                                                                   // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [15:0] rsp_xbar_demux_001_src1_channel;                                                                                // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                                  // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_001_src2_endofpacket;                                                                            // rsp_xbar_demux_001:src2_endofpacket -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_001_src2_valid;                                                                                  // rsp_xbar_demux_001:src2_valid -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_001_src2_startofpacket;                                                                          // rsp_xbar_demux_001:src2_startofpacket -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src2_data;                                                                                   // rsp_xbar_demux_001:src2_data -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_demux_001_src2_channel;                                                                                // rsp_xbar_demux_001:src2_channel -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_001_src3_endofpacket;                                                                            // rsp_xbar_demux_001:src3_endofpacket -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_001_src3_valid;                                                                                  // rsp_xbar_demux_001:src3_valid -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_001_src3_startofpacket;                                                                          // rsp_xbar_demux_001:src3_startofpacket -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src3_data;                                                                                   // rsp_xbar_demux_001:src3_data -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_demux_001_src3_channel;                                                                                // rsp_xbar_demux_001:src3_channel -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                            // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                  // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                          // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_002_src0_data;                                                                                   // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [15:0] rsp_xbar_demux_002_src0_channel;                                                                                // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                  // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                            // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                                  // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                          // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_002_src1_data;                                                                                   // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [15:0] rsp_xbar_demux_002_src1_channel;                                                                                // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                                  // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                            // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                  // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                          // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src0_data;                                                                                   // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [15:0] rsp_xbar_demux_003_src0_channel;                                                                                // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                  // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                            // rsp_xbar_demux_003:src1_endofpacket -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                                  // rsp_xbar_demux_003:src1_valid -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                                          // rsp_xbar_demux_003:src1_startofpacket -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src1_data;                                                                                   // rsp_xbar_demux_003:src1_data -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_demux_003_src1_channel;                                                                                // rsp_xbar_demux_003:src1_channel -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_003_src2_endofpacket;                                                                            // rsp_xbar_demux_003:src2_endofpacket -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_003_src2_valid;                                                                                  // rsp_xbar_demux_003:src2_valid -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_003_src2_startofpacket;                                                                          // rsp_xbar_demux_003:src2_startofpacket -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src2_data;                                                                                   // rsp_xbar_demux_003:src2_data -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_demux_003_src2_channel;                                                                                // rsp_xbar_demux_003:src2_channel -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_003_src3_endofpacket;                                                                            // rsp_xbar_demux_003:src3_endofpacket -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_003_src3_valid;                                                                                  // rsp_xbar_demux_003:src3_valid -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_003_src3_startofpacket;                                                                          // rsp_xbar_demux_003:src3_startofpacket -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src3_data;                                                                                   // rsp_xbar_demux_003:src3_data -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_demux_003_src3_channel;                                                                                // rsp_xbar_demux_003:src3_channel -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_003_src4_endofpacket;                                                                            // rsp_xbar_demux_003:src4_endofpacket -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_003_src4_valid;                                                                                  // rsp_xbar_demux_003:src4_valid -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_003_src4_startofpacket;                                                                          // rsp_xbar_demux_003:src4_startofpacket -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src4_data;                                                                                   // rsp_xbar_demux_003:src4_data -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_demux_003_src4_channel;                                                                                // rsp_xbar_demux_003:src4_channel -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                            // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                  // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                          // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_004_src0_data;                                                                                   // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [15:0] rsp_xbar_demux_004_src0_channel;                                                                                // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                  // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                            // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                  // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                          // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_005_src0_data;                                                                                   // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [15:0] rsp_xbar_demux_005_src0_channel;                                                                                // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                                  // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                            // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                                  // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                          // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [106:0] rsp_xbar_demux_006_src0_data;                                                                                   // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [15:0] rsp_xbar_demux_006_src0_channel;                                                                                // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                                  // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                            // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                                  // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                          // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [106:0] rsp_xbar_demux_007_src0_data;                                                                                   // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [15:0] rsp_xbar_demux_007_src0_channel;                                                                                // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                                  // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                            // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                                  // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                          // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [106:0] rsp_xbar_demux_008_src0_data;                                                                                   // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [15:0] rsp_xbar_demux_008_src0_channel;                                                                                // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                                  // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                            // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                                  // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                          // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [106:0] rsp_xbar_demux_009_src0_data;                                                                                   // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [15:0] rsp_xbar_demux_009_src0_channel;                                                                                // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                                  // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_009_src1_endofpacket;                                                                            // rsp_xbar_demux_009:src1_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire          rsp_xbar_demux_009_src1_valid;                                                                                  // rsp_xbar_demux_009:src1_valid -> rsp_xbar_mux_002:sink0_valid
	wire          rsp_xbar_demux_009_src1_startofpacket;                                                                          // rsp_xbar_demux_009:src1_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_009_src1_data;                                                                                   // rsp_xbar_demux_009:src1_data -> rsp_xbar_mux_002:sink0_data
	wire   [15:0] rsp_xbar_demux_009_src1_channel;                                                                                // rsp_xbar_demux_009:src1_channel -> rsp_xbar_mux_002:sink0_channel
	wire          rsp_xbar_demux_009_src1_ready;                                                                                  // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_009:src1_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                            // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                                  // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                          // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [106:0] rsp_xbar_demux_010_src0_data;                                                                                   // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [15:0] rsp_xbar_demux_010_src0_channel;                                                                                // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                                  // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_010_src1_endofpacket;                                                                            // rsp_xbar_demux_010:src1_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire          rsp_xbar_demux_010_src1_valid;                                                                                  // rsp_xbar_demux_010:src1_valid -> rsp_xbar_mux_002:sink1_valid
	wire          rsp_xbar_demux_010_src1_startofpacket;                                                                          // rsp_xbar_demux_010:src1_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_010_src1_data;                                                                                   // rsp_xbar_demux_010:src1_data -> rsp_xbar_mux_002:sink1_data
	wire   [15:0] rsp_xbar_demux_010_src1_channel;                                                                                // rsp_xbar_demux_010:src1_channel -> rsp_xbar_mux_002:sink1_channel
	wire          rsp_xbar_demux_010_src1_ready;                                                                                  // rsp_xbar_mux_002:sink1_ready -> rsp_xbar_demux_010:src1_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                            // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                                  // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                          // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [106:0] rsp_xbar_demux_011_src0_data;                                                                                   // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire   [15:0] rsp_xbar_demux_011_src0_channel;                                                                                // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                                  // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                            // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                                  // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_002:sink2_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                          // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_012_src0_data;                                                                                   // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_002:sink2_data
	wire   [15:0] rsp_xbar_demux_012_src0_channel;                                                                                // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_002:sink2_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                                  // rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                            // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                                  // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_002:sink3_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                          // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_013_src0_data;                                                                                   // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_002:sink3_data
	wire   [15:0] rsp_xbar_demux_013_src0_channel;                                                                                // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_002:sink3_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                                  // rsp_xbar_mux_002:sink3_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_013_src1_endofpacket;                                                                            // rsp_xbar_demux_013:src1_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire          rsp_xbar_demux_013_src1_valid;                                                                                  // rsp_xbar_demux_013:src1_valid -> rsp_xbar_mux_003:sink0_valid
	wire          rsp_xbar_demux_013_src1_startofpacket;                                                                          // rsp_xbar_demux_013:src1_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_013_src1_data;                                                                                   // rsp_xbar_demux_013:src1_data -> rsp_xbar_mux_003:sink0_data
	wire   [15:0] rsp_xbar_demux_013_src1_channel;                                                                                // rsp_xbar_demux_013:src1_channel -> rsp_xbar_mux_003:sink0_channel
	wire          rsp_xbar_demux_013_src1_ready;                                                                                  // rsp_xbar_mux_003:sink0_ready -> rsp_xbar_demux_013:src1_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                            // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_002:sink4_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                                  // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_002:sink4_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                          // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_002:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_014_src0_data;                                                                                   // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_002:sink4_data
	wire   [15:0] rsp_xbar_demux_014_src0_channel;                                                                                // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_002:sink4_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                                  // rsp_xbar_mux_002:sink4_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_014_src1_endofpacket;                                                                            // rsp_xbar_demux_014:src1_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire          rsp_xbar_demux_014_src1_valid;                                                                                  // rsp_xbar_demux_014:src1_valid -> rsp_xbar_mux_003:sink1_valid
	wire          rsp_xbar_demux_014_src1_startofpacket;                                                                          // rsp_xbar_demux_014:src1_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_014_src1_data;                                                                                   // rsp_xbar_demux_014:src1_data -> rsp_xbar_mux_003:sink1_data
	wire   [15:0] rsp_xbar_demux_014_src1_channel;                                                                                // rsp_xbar_demux_014:src1_channel -> rsp_xbar_mux_003:sink1_channel
	wire          rsp_xbar_demux_014_src1_ready;                                                                                  // rsp_xbar_mux_003:sink1_ready -> rsp_xbar_demux_014:src1_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                            // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_002:sink5_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                                  // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_002:sink5_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                          // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_002:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_015_src0_data;                                                                                   // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_002:sink5_data
	wire   [15:0] rsp_xbar_demux_015_src0_channel;                                                                                // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_002:sink5_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                                  // rsp_xbar_mux_002:sink5_ready -> rsp_xbar_demux_015:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                                    // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                                  // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [106:0] limiter_cmd_src_data;                                                                                           // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [15:0] limiter_cmd_src_channel;                                                                                        // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                          // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                   // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                         // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                                 // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_src_data;                                                                                          // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [15:0] rsp_xbar_mux_src_channel;                                                                                       // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                         // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                                // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                      // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                              // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [106:0] addr_router_001_src_data;                                                                                       // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [15:0] addr_router_001_src_channel;                                                                                    // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                                      // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                               // rsp_xbar_mux_001:src_endofpacket -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                     // rsp_xbar_mux_001:src_valid -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                             // rsp_xbar_mux_001:src_startofpacket -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_mux_001_src_data;                                                                                      // rsp_xbar_mux_001:src_data -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_mux_001_src_channel;                                                                                   // rsp_xbar_mux_001:src_channel -> nios2_communication_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                     // nios2_communication_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                                // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                      // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                              // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [106:0] addr_router_002_src_data;                                                                                       // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [15:0] addr_router_002_src_channel;                                                                                    // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                                      // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_mux_002_src_endofpacket;                                                                               // rsp_xbar_mux_002:src_endofpacket -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_002_src_valid;                                                                                     // rsp_xbar_mux_002:src_valid -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_002_src_startofpacket;                                                                             // rsp_xbar_mux_002:src_startofpacket -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_mux_002_src_data;                                                                                      // rsp_xbar_mux_002:src_data -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_mux_002_src_channel;                                                                                   // rsp_xbar_mux_002:src_channel -> nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_002_src_ready;                                                                                     // nios2_car_controll_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_002:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                                // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                              // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [106:0] limiter_001_cmd_src_data;                                                                                       // limiter_001:cmd_src_data -> cmd_xbar_demux_003:sink_data
	wire   [15:0] limiter_001_cmd_src_channel;                                                                                    // limiter_001:cmd_src_channel -> cmd_xbar_demux_003:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                                      // cmd_xbar_demux_003:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_003_src_endofpacket;                                                                               // rsp_xbar_mux_003:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_003_src_valid;                                                                                     // rsp_xbar_mux_003:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_003_src_startofpacket;                                                                             // rsp_xbar_mux_003:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_003_src_data;                                                                                      // rsp_xbar_mux_003:src_data -> limiter_001:rsp_sink_data
	wire   [15:0] rsp_xbar_mux_003_src_channel;                                                                                   // rsp_xbar_mux_003:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_003_src_ready;                                                                                     // limiter_001:rsp_sink_ready -> rsp_xbar_mux_003:src_ready
	wire          addr_router_004_src_endofpacket;                                                                                // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          addr_router_004_src_valid;                                                                                      // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire          addr_router_004_src_startofpacket;                                                                              // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [106:0] addr_router_004_src_data;                                                                                       // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire   [15:0] addr_router_004_src_channel;                                                                                    // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire          addr_router_004_src_ready;                                                                                      // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire          rsp_xbar_demux_003_src1_ready;                                                                                  // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_003:src1_ready
	wire          addr_router_005_src_endofpacket;                                                                                // addr_router_005:src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          addr_router_005_src_valid;                                                                                      // addr_router_005:src_valid -> cmd_xbar_demux_005:sink_valid
	wire          addr_router_005_src_startofpacket;                                                                              // addr_router_005:src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire  [106:0] addr_router_005_src_data;                                                                                       // addr_router_005:src_data -> cmd_xbar_demux_005:sink_data
	wire   [15:0] addr_router_005_src_channel;                                                                                    // addr_router_005:src_channel -> cmd_xbar_demux_005:sink_channel
	wire          addr_router_005_src_ready;                                                                                      // cmd_xbar_demux_005:sink_ready -> addr_router_005:src_ready
	wire          rsp_xbar_demux_003_src2_ready;                                                                                  // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_003:src2_ready
	wire          addr_router_006_src_endofpacket;                                                                                // addr_router_006:src_endofpacket -> cmd_xbar_demux_006:sink_endofpacket
	wire          addr_router_006_src_valid;                                                                                      // addr_router_006:src_valid -> cmd_xbar_demux_006:sink_valid
	wire          addr_router_006_src_startofpacket;                                                                              // addr_router_006:src_startofpacket -> cmd_xbar_demux_006:sink_startofpacket
	wire  [106:0] addr_router_006_src_data;                                                                                       // addr_router_006:src_data -> cmd_xbar_demux_006:sink_data
	wire   [15:0] addr_router_006_src_channel;                                                                                    // addr_router_006:src_channel -> cmd_xbar_demux_006:sink_channel
	wire          addr_router_006_src_ready;                                                                                      // cmd_xbar_demux_006:sink_ready -> addr_router_006:src_ready
	wire          rsp_xbar_demux_003_src3_ready;                                                                                  // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_003:src3_ready
	wire          addr_router_007_src_endofpacket;                                                                                // addr_router_007:src_endofpacket -> cmd_xbar_demux_007:sink_endofpacket
	wire          addr_router_007_src_valid;                                                                                      // addr_router_007:src_valid -> cmd_xbar_demux_007:sink_valid
	wire          addr_router_007_src_startofpacket;                                                                              // addr_router_007:src_startofpacket -> cmd_xbar_demux_007:sink_startofpacket
	wire  [106:0] addr_router_007_src_data;                                                                                       // addr_router_007:src_data -> cmd_xbar_demux_007:sink_data
	wire   [15:0] addr_router_007_src_channel;                                                                                    // addr_router_007:src_channel -> cmd_xbar_demux_007:sink_channel
	wire          addr_router_007_src_ready;                                                                                      // cmd_xbar_demux_007:sink_ready -> addr_router_007:src_ready
	wire          rsp_xbar_demux_003_src4_ready;                                                                                  // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_003:src4_ready
	wire          addr_router_008_src_endofpacket;                                                                                // addr_router_008:src_endofpacket -> cmd_xbar_demux_008:sink_endofpacket
	wire          addr_router_008_src_valid;                                                                                      // addr_router_008:src_valid -> cmd_xbar_demux_008:sink_valid
	wire          addr_router_008_src_startofpacket;                                                                              // addr_router_008:src_startofpacket -> cmd_xbar_demux_008:sink_startofpacket
	wire  [106:0] addr_router_008_src_data;                                                                                       // addr_router_008:src_data -> cmd_xbar_demux_008:sink_data
	wire   [15:0] addr_router_008_src_channel;                                                                                    // addr_router_008:src_channel -> cmd_xbar_demux_008:sink_channel
	wire          addr_router_008_src_ready;                                                                                      // cmd_xbar_demux_008:sink_ready -> addr_router_008:src_ready
	wire          rsp_xbar_demux_001_src2_ready;                                                                                  // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_001:src2_ready
	wire          addr_router_009_src_endofpacket;                                                                                // addr_router_009:src_endofpacket -> cmd_xbar_demux_009:sink_endofpacket
	wire          addr_router_009_src_valid;                                                                                      // addr_router_009:src_valid -> cmd_xbar_demux_009:sink_valid
	wire          addr_router_009_src_startofpacket;                                                                              // addr_router_009:src_startofpacket -> cmd_xbar_demux_009:sink_startofpacket
	wire  [106:0] addr_router_009_src_data;                                                                                       // addr_router_009:src_data -> cmd_xbar_demux_009:sink_data
	wire   [15:0] addr_router_009_src_channel;                                                                                    // addr_router_009:src_channel -> cmd_xbar_demux_009:sink_channel
	wire          addr_router_009_src_ready;                                                                                      // cmd_xbar_demux_009:sink_ready -> addr_router_009:src_ready
	wire          rsp_xbar_demux_001_src3_ready;                                                                                  // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_001:src3_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                                   // cmd_xbar_mux:src_endofpacket -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                         // cmd_xbar_mux:src_valid -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                                 // cmd_xbar_mux:src_startofpacket -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_src_data;                                                                                          // cmd_xbar_mux:src_data -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_src_channel;                                                                                       // cmd_xbar_mux:src_channel -> nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                         // nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                      // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                            // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                    // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [106:0] id_router_src_data;                                                                                             // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [15:0] id_router_src_channel;                                                                                          // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                            // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                               // cmd_xbar_mux_001:src_endofpacket -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                     // cmd_xbar_mux_001:src_valid -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                             // cmd_xbar_mux_001:src_startofpacket -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_001_src_data;                                                                                      // cmd_xbar_mux_001:src_data -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_001_src_channel;                                                                                   // cmd_xbar_mux_001:src_channel -> main_memory_communication_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                     // main_memory_communication_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                                  // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                        // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                                // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [106:0] id_router_001_src_data;                                                                                         // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [15:0] id_router_001_src_channel;                                                                                      // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                        // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                               // cmd_xbar_mux_002:src_endofpacket -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                                     // cmd_xbar_mux_002:src_valid -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                             // cmd_xbar_mux_002:src_startofpacket -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_002_src_data;                                                                                      // cmd_xbar_mux_002:src_data -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_002_src_channel;                                                                                   // cmd_xbar_mux_002:src_channel -> sdram_communication_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                                     // sdram_communication_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                                  // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                        // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                                // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [106:0] id_router_002_src_data;                                                                                         // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [15:0] id_router_002_src_channel;                                                                                      // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                        // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                               // cmd_xbar_mux_003:src_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                                     // cmd_xbar_mux_003:src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                             // cmd_xbar_mux_003:src_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_003_src_data;                                                                                      // cmd_xbar_mux_003:src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_003_src_channel;                                                                                   // cmd_xbar_mux_003:src_channel -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                                     // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                                  // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                        // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                                // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [106:0] id_router_003_src_data;                                                                                         // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [15:0] id_router_003_src_channel;                                                                                      // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                        // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                                  // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                                  // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                        // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                                // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [106:0] id_router_004_src_data;                                                                                         // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [15:0] id_router_004_src_channel;                                                                                      // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                        // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                                  // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                                  // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                        // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                                // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [106:0] id_router_005_src_data;                                                                                         // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [15:0] id_router_005_src_channel;                                                                                      // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                        // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                                  // tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                                  // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                        // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                                // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [106:0] id_router_006_src_data;                                                                                         // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [15:0] id_router_006_src_channel;                                                                                      // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                        // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                                  // jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                                  // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                        // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                                // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [106:0] id_router_007_src_data;                                                                                         // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [15:0] id_router_007_src_channel;                                                                                      // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                        // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                                  // shared_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_008_src_endofpacket;                                                                                  // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                        // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                                // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [106:0] id_router_008_src_data;                                                                                         // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [15:0] id_router_008_src_channel;                                                                                      // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                        // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_mux_009_src_endofpacket;                                                                               // cmd_xbar_mux_009:src_endofpacket -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_009_src_valid;                                                                                     // cmd_xbar_mux_009:src_valid -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_009_src_startofpacket;                                                                             // cmd_xbar_mux_009:src_startofpacket -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_009_src_data;                                                                                      // cmd_xbar_mux_009:src_data -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_009_src_channel;                                                                                   // cmd_xbar_mux_009:src_channel -> mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_009_src_ready;                                                                                     // mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	wire          id_router_009_src_endofpacket;                                                                                  // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                        // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                                // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [106:0] id_router_009_src_data;                                                                                         // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [15:0] id_router_009_src_channel;                                                                                      // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                        // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_mux_010_src_endofpacket;                                                                               // cmd_xbar_mux_010:src_endofpacket -> interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_010_src_valid;                                                                                     // cmd_xbar_mux_010:src_valid -> interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_010_src_startofpacket;                                                                             // cmd_xbar_mux_010:src_startofpacket -> interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_010_src_data;                                                                                      // cmd_xbar_mux_010:src_data -> interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_010_src_channel;                                                                                   // cmd_xbar_mux_010:src_channel -> interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_010_src_ready;                                                                                     // interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_010:src_ready
	wire          id_router_010_src_endofpacket;                                                                                  // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                        // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                                // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [106:0] id_router_010_src_data;                                                                                         // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [15:0] id_router_010_src_channel;                                                                                      // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                        // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_001_src11_ready;                                                                                 // pio_communication_led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire          id_router_011_src_endofpacket;                                                                                  // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                        // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                                // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [106:0] id_router_011_src_data;                                                                                         // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [15:0] id_router_011_src_channel;                                                                                      // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                        // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_002_src2_ready;                                                                                  // shared_memory_s2_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src2_ready
	wire          id_router_012_src_endofpacket;                                                                                  // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                        // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                                // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [106:0] id_router_012_src_data;                                                                                         // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [15:0] id_router_012_src_channel;                                                                                      // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                        // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_mux_013_src_endofpacket;                                                                               // cmd_xbar_mux_013:src_endofpacket -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_013_src_valid;                                                                                     // cmd_xbar_mux_013:src_valid -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_013_src_startofpacket;                                                                             // cmd_xbar_mux_013:src_startofpacket -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_013_src_data;                                                                                      // cmd_xbar_mux_013:src_data -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_013_src_channel;                                                                                   // cmd_xbar_mux_013:src_channel -> main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_013_src_ready;                                                                                     // main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_013:src_ready
	wire          id_router_013_src_endofpacket;                                                                                  // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                        // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                                // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [106:0] id_router_013_src_data;                                                                                         // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [15:0] id_router_013_src_channel;                                                                                      // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                        // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_mux_014_src_endofpacket;                                                                               // cmd_xbar_mux_014:src_endofpacket -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_014_src_valid;                                                                                     // cmd_xbar_mux_014:src_valid -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_014_src_startofpacket;                                                                             // cmd_xbar_mux_014:src_startofpacket -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_014_src_data;                                                                                      // cmd_xbar_mux_014:src_data -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_014_src_channel;                                                                                   // cmd_xbar_mux_014:src_channel -> nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_014_src_ready;                                                                                     // nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_014:src_ready
	wire          id_router_014_src_endofpacket;                                                                                  // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                        // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                                // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [106:0] id_router_014_src_data;                                                                                         // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [15:0] id_router_014_src_channel;                                                                                      // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                        // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_002_src5_ready;                                                                                  // jtag_uart_carControl_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_002:src5_ready
	wire          id_router_015_src_endofpacket;                                                                                  // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                        // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                                // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [106:0] id_router_015_src_data;                                                                                         // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [15:0] id_router_015_src_channel;                                                                                      // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                        // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire   [15:0] limiter_cmd_valid_data;                                                                                         // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [15:0] limiter_001_cmd_valid_data;                                                                                     // limiter_001:cmd_src_valid -> cmd_xbar_demux_003:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                                       // jtag_uart_communication:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                       // sgdma_rx:csr_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                       // sgdma_tx:csr_irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                                       // interval_timer:irq -> irq_mapper:receiver3_irq
	wire   [31:0] nios2_communication_d_irq_irq;                                                                                  // irq_mapper:sender_irq -> nios2_communication:d_irq
	wire          irq_mapper_001_receiver0_irq;                                                                                   // jtag_uart_carControl:av_irq -> irq_mapper_001:receiver0_irq
	wire   [31:0] nios2_car_controll_d_irq_irq;                                                                                   // irq_mapper_001:sender_irq -> nios2_car_controll:d_irq

	nios_system_nios2_communication nios2_communication (
		.clk                                   (clk_clk),                                                                            //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                                    //                   reset_n.reset_n
		.d_address                             (nios2_communication_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_communication_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_communication_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_communication_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_communication_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_communication_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_communication_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_communication_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_communication_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_communication_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_communication_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_communication_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (nios2_communication_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (nios2_communication_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_communication_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                                    // custom_instruction_master.readra
	);

	nios_system_main_memory_communication main_memory_communication (
		.clk        (clk_clk),                                                                //   clk1.clk
		.address    (main_memory_communication_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (main_memory_communication_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (main_memory_communication_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (main_memory_communication_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (main_memory_communication_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (main_memory_communication_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (main_memory_communication_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                                          // reset1.reset
	);

	nios_system_jtag_uart_communication jtag_uart_communication (
		.clk            (clk_clk),                                                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                              //               irq.irq
	);

	nios_system_tse_mac tse_mac (
		.ff_tx_data  (sgdma_tx_out_data),                                               //                      transmit.data
		.ff_tx_eop   (sgdma_tx_out_endofpacket),                                        //                              .endofpacket
		.ff_tx_err   (sgdma_tx_out_error),                                              //                              .error
		.ff_tx_mod   (sgdma_tx_out_empty),                                              //                              .empty
		.ff_tx_rdy   (sgdma_tx_out_ready),                                              //                              .ready
		.ff_tx_sop   (sgdma_tx_out_startofpacket),                                      //                              .startofpacket
		.ff_tx_wren  (sgdma_tx_out_valid),                                              //                              .valid
		.ff_tx_clk   (clk_clk),                                                         //      receive_clock_connection.clk
		.ff_rx_data  (tse_mac_receive_data),                                            //                       receive.data
		.ff_rx_dval  (tse_mac_receive_valid),                                           //                              .valid
		.ff_rx_eop   (tse_mac_receive_endofpacket),                                     //                              .endofpacket
		.ff_rx_mod   (tse_mac_receive_empty),                                           //                              .empty
		.ff_rx_rdy   (tse_mac_receive_ready),                                           //                              .ready
		.ff_rx_sop   (tse_mac_receive_startofpacket),                                   //                              .startofpacket
		.rx_err      (tse_mac_receive_error),                                           //                              .error
		.ff_rx_clk   (clk_clk),                                                         //     transmit_clock_connection.clk
		.address     (tse_mac_control_port_translator_avalon_anti_slave_0_address),     //                  control_port.address
		.readdata    (tse_mac_control_port_translator_avalon_anti_slave_0_readdata),    //                              .readdata
		.read        (tse_mac_control_port_translator_avalon_anti_slave_0_read),        //                              .read
		.writedata   (tse_mac_control_port_translator_avalon_anti_slave_0_writedata),   //                              .writedata
		.write       (tse_mac_control_port_translator_avalon_anti_slave_0_write),       //                              .write
		.waitrequest (tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest), //                              .waitrequest
		.clk         (clk_clk),                                                         // control_port_clock_connection.clk
		.reset       (rst_controller_reset_out_reset),                                  //              reset_connection.reset
		.rgmii_in    (tse_mac_conduit_connection_rgmii_in),                             //            conduit_connection.export
		.rgmii_out   (tse_mac_conduit_connection_rgmii_out),                            //                              .export
		.rx_control  (tse_mac_conduit_connection_rx_control),                           //                              .export
		.tx_control  (tse_mac_conduit_connection_tx_control),                           //                              .export
		.tx_clk      (tse_mac_conduit_connection_tx_clk),                               //                              .export
		.rx_clk      (tse_mac_conduit_connection_rx_clk),                               //                              .export
		.set_10      (tse_mac_conduit_connection_set_10),                               //                              .export
		.set_1000    (tse_mac_conduit_connection_set_1000),                             //                              .export
		.ena_10      (tse_mac_conduit_connection_ena_10),                               //                              .export
		.eth_mode    (tse_mac_conduit_connection_eth_mode),                             //                              .export
		.mdio_out    (tse_mac_conduit_connection_mdio_out),                             //                              .export
		.mdio_oen    (tse_mac_conduit_connection_mdio_oen),                             //                              .export
		.mdio_in     (tse_mac_conduit_connection_mdio_in),                              //                              .export
		.mdc         (tse_mac_conduit_connection_mdc)                                   //                              .export
	);

	nios_system_sgdma_rx sgdma_rx (
		.clk                           (clk_clk),                                                //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),                        //            reset.reset_n
		.csr_chipselect                (sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (sgdma_rx_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (sgdma_rx_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (sgdma_rx_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (sgdma_rx_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (sgdma_rx_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (sgdma_rx_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (sgdma_rx_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_rx_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (sgdma_rx_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (irq_mapper_receiver1_irq),                               //          csr_irq.irq
		.m_write_waitrequest           (sgdma_rx_m_write_waitrequest),                           //          m_write.waitrequest
		.m_write_address               (sgdma_rx_m_write_address),                               //                 .address
		.m_write_write                 (sgdma_rx_m_write_write),                                 //                 .write
		.m_write_writedata             (sgdma_rx_m_write_writedata),                             //                 .writedata
		.m_write_byteenable            (sgdma_rx_m_write_byteenable),                            //                 .byteenable
		.in_startofpacket              (tse_mac_receive_startofpacket),                          //               in.startofpacket
		.in_endofpacket                (tse_mac_receive_endofpacket),                            //                 .endofpacket
		.in_empty                      (tse_mac_receive_empty),                                  //                 .empty
		.in_data                       (tse_mac_receive_data),                                   //                 .data
		.in_valid                      (tse_mac_receive_valid),                                  //                 .valid
		.in_ready                      (tse_mac_receive_ready),                                  //                 .ready
		.in_error                      (tse_mac_receive_error)                                   //                 .error
	);

	nios_system_sgdma_tx sgdma_tx (
		.clk                           (clk_clk),                                                //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),                        //            reset.reset_n
		.csr_chipselect                (sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (sgdma_tx_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (sgdma_tx_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (sgdma_tx_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (sgdma_tx_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (sgdma_tx_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (sgdma_tx_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (sgdma_tx_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_tx_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (sgdma_tx_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (irq_mapper_receiver2_irq),                               //          csr_irq.irq
		.m_read_readdata               (sgdma_tx_m_read_readdata),                               //           m_read.readdata
		.m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),                          //                 .readdatavalid
		.m_read_waitrequest            (sgdma_tx_m_read_waitrequest),                            //                 .waitrequest
		.m_read_address                (sgdma_tx_m_read_address),                                //                 .address
		.m_read_read                   (sgdma_tx_m_read_read),                                   //                 .read
		.out_data                      (sgdma_tx_out_data),                                      //              out.data
		.out_valid                     (sgdma_tx_out_valid),                                     //                 .valid
		.out_ready                     (sgdma_tx_out_ready),                                     //                 .ready
		.out_endofpacket               (sgdma_tx_out_endofpacket),                               //                 .endofpacket
		.out_startofpacket             (sgdma_tx_out_startofpacket),                             //                 .startofpacket
		.out_empty                     (sgdma_tx_out_empty),                                     //                 .empty
		.out_error                     (sgdma_tx_out_error)                                      //                 .error
	);

	nios_system_descriptor_memory descriptor_memory (
		.clk        (clk_clk),                                                        //   clk1.clk
		.address    (descriptor_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (descriptor_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (descriptor_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (descriptor_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (descriptor_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                                  // reset1.reset
	);

	nios_system_nios2_car_controll nios2_car_controll (
		.clk                                   (clk_clk),                                                                           //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                                   //                   reset_n.reset_n
		.d_address                             (nios2_car_controll_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_car_controll_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_car_controll_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_car_controll_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_car_controll_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_car_controll_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_car_controll_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_car_controll_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_car_controll_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_car_controll_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_car_controll_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_car_controll_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (nios2_car_controll_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (nios2_car_controll_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_car_controll_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                                   // custom_instruction_master.readra
	);

	nios_system_shared_memory shared_memory (
		.clk         (clk_clk),                                                    //   clk1.clk
		.address     (shared_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect  (shared_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken       (shared_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata    (shared_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write       (shared_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata   (shared_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable  (shared_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                             // reset1.reset
		.address2    (shared_memory_s2_translator_avalon_anti_slave_0_address),    //     s2.address
		.chipselect2 (shared_memory_s2_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken2      (shared_memory_s2_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata2   (shared_memory_s2_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write2      (shared_memory_s2_translator_avalon_anti_slave_0_write),      //       .write
		.writedata2  (shared_memory_s2_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable2 (shared_memory_s2_translator_avalon_anti_slave_0_byteenable)  //       .byteenable
	);

	nios_system_main_memory_car_controll main_memory_car_controll (
		.clk        (clk_clk),                                                               //   clk1.clk
		.address    (main_memory_car_controll_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (main_memory_car_controll_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (main_memory_car_controll_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (main_memory_car_controll_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (main_memory_car_controll_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (main_memory_car_controll_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (main_memory_car_controll_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                                         // reset1.reset
	);

	nios_system_mutex_shared_memory mutex_shared_memory (
		.clk           (clk_clk),                                                          //   clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                  // reset.reset_n
		.address       (mutex_shared_memory_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.chipselect    (mutex_shared_memory_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.data_from_cpu (mutex_shared_memory_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.data_to_cpu   (mutex_shared_memory_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.read          (mutex_shared_memory_s1_translator_avalon_anti_slave_0_read),       //      .read
		.write         (mutex_shared_memory_s1_translator_avalon_anti_slave_0_write)       //      .write
	);

	nios_system_jtag_uart_communication jtag_uart_carcontrol (
		.clk            (clk_clk),                                                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                                   //             reset.reset_n
		.av_chipselect  (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver0_irq)                                                       //               irq.irq
	);

	nios_system_interval_timer interval_timer (
		.clk        (clk_clk),                                                     //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                             // reset.reset_n
		.address    (interval_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (interval_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (interval_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (interval_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~interval_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                                     //   irq.irq
	);

	nios_system_pio_communication_led pio_communication_led (
		.clk        (clk_clk),                                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                                    //               reset.reset_n
		.address    (pio_communication_led_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_communication_led_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_communication_led_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_communication_led_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_communication_led_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (pio_communication_led_external_connection_export)                    // external_connection.export
	);

	nios_system_sdram_communication sdram_communication (
		.clk            (clk_clk),                                                             //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                                 // reset.reset_n
		.az_addr        (sdram_communication_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_communication_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_communication_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_communication_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_communication_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_communication_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_communication_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_communication_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_communication_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_communication_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_communication_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_communication_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_communication_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_communication_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_communication_wire_dq),                                         //      .export
		.zs_dqm         (sdram_communication_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_communication_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_communication_wire_we_n)                                        //      .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_communication_instruction_master_translator (
		.clk                   (clk_clk),                                                                                   //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                            //                     reset.reset
		.uav_address           (nios2_communication_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_communication_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_communication_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_communication_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_communication_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_communication_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_communication_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_communication_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_communication_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_communication_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_communication_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_communication_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_communication_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (nios2_communication_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_communication_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_communication_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                                      //               (terminated)
		.av_byteenable         (4'b1111),                                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                                      //               (terminated)
		.av_write              (1'b0),                                                                                      //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                                      //               (terminated)
		.av_lock               (1'b0),                                                                                      //               (terminated)
		.av_debugaccess        (1'b0),                                                                                      //               (terminated)
		.uav_clken             (),                                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_communication_data_master_translator (
		.clk                   (clk_clk),                                                                            //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address           (nios2_communication_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_communication_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_communication_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_communication_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_communication_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_communication_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_communication_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_communication_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_communication_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_communication_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_communication_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_communication_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_communication_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (nios2_communication_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_communication_data_master_read),                                               //                          .read
		.av_readdata           (nios2_communication_data_master_readdata),                                           //                          .readdata
		.av_write              (nios2_communication_data_master_write),                                              //                          .write
		.av_writedata          (nios2_communication_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_communication_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                                               //               (terminated)
		.av_readdatavalid      (),                                                                                   //               (terminated)
		.av_lock               (1'b0),                                                                               //               (terminated)
		.uav_clken             (),                                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_car_controll_data_master_translator (
		.clk                   (clk_clk),                                                                           //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                    //                     reset.reset
		.uav_address           (nios2_car_controll_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_car_controll_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_car_controll_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_car_controll_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_car_controll_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_car_controll_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_car_controll_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_car_controll_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_car_controll_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_car_controll_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_car_controll_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_car_controll_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_car_controll_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (nios2_car_controll_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_car_controll_data_master_read),                                               //                          .read
		.av_readdata           (nios2_car_controll_data_master_readdata),                                           //                          .readdata
		.av_write              (nios2_car_controll_data_master_write),                                              //                          .write
		.av_writedata          (nios2_car_controll_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_car_controll_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                              //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                              //               (terminated)
		.av_begintransfer      (1'b0),                                                                              //               (terminated)
		.av_chipselect         (1'b0),                                                                              //               (terminated)
		.av_readdatavalid      (),                                                                                  //               (terminated)
		.av_lock               (1'b0),                                                                              //               (terminated)
		.uav_clken             (),                                                                                  //               (terminated)
		.av_clken              (1'b1)                                                                               //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (19),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_car_controll_instruction_master_translator (
		.clk                   (clk_clk),                                                                                  //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                           //                     reset.reset
		.uav_address           (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_car_controll_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_car_controll_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (nios2_car_controll_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_car_controll_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_car_controll_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                                     //               (terminated)
		.av_byteenable         (4'b1111),                                                                                  //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                     //               (terminated)
		.av_begintransfer      (1'b0),                                                                                     //               (terminated)
		.av_chipselect         (1'b0),                                                                                     //               (terminated)
		.av_write              (1'b0),                                                                                     //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                                     //               (terminated)
		.av_lock               (1'b0),                                                                                     //               (terminated)
		.av_debugaccess        (1'b0),                                                                                     //               (terminated)
		.uav_clken             (),                                                                                         //               (terminated)
		.av_clken              (1'b1)                                                                                      //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_m_write_translator (
		.clk                   (clk_clk),                                                             //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                     reset.reset
		.uav_address           (sgdma_rx_m_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_m_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_m_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_m_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_m_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_m_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_m_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_m_write_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (sgdma_rx_m_write_byteenable),                                         //                          .byteenable
		.av_write              (sgdma_rx_m_write_write),                                              //                          .write
		.av_writedata          (sgdma_rx_m_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                //               (terminated)
		.av_begintransfer      (1'b0),                                                                //               (terminated)
		.av_chipselect         (1'b0),                                                                //               (terminated)
		.av_read               (1'b0),                                                                //               (terminated)
		.av_readdata           (),                                                                    //               (terminated)
		.av_readdatavalid      (),                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                //               (terminated)
		.av_debugaccess        (1'b0),                                                                //               (terminated)
		.uav_clken             (),                                                                    //               (terminated)
		.av_clken              (1'b1)                                                                 //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_m_read_translator (
		.clk                   (clk_clk),                                                            //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address           (sgdma_tx_m_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_m_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_m_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_m_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_m_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_m_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_m_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_m_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_tx_m_read_read),                                               //                          .read
		.av_readdata           (sgdma_tx_m_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_tx_m_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_byteenable         (4'b1111),                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_write              (1'b0),                                                               //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                               //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_descriptor_read_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_rx_descriptor_read_read),                                               //                          .read
		.av_readdata           (sgdma_rx_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_rx_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_descriptor_write_translator (
		.clk                   (clk_clk),                                                                      //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                     reset.reset
		.uav_address           (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write              (sgdma_rx_descriptor_write_write),                                              //                          .write
		.av_writedata          (sgdma_rx_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                         //               (terminated)
		.av_byteenable         (4'b1111),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_read               (1'b0),                                                                         //               (terminated)
		.av_readdata           (),                                                                             //               (terminated)
		.av_readdatavalid      (),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.av_debugaccess        (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_descriptor_read_translator (
		.clk                   (clk_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_tx_descriptor_read_read),                                               //                          .read
		.av_readdata           (sgdma_tx_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_tx_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_descriptor_write_translator (
		.clk                   (clk_clk),                                                                      //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                     reset.reset
		.uav_address           (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write              (sgdma_tx_descriptor_write_write),                                              //                          .write
		.av_writedata          (sgdma_tx_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                         //               (terminated)
		.av_byteenable         (4'b1111),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_read               (1'b0),                                                                         //               (terminated)
		.av_readdata           (),                                                                             //               (terminated)
		.av_readdatavalid      (),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.av_debugaccess        (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_communication_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                   //                    reset.reset
		.uav_address           (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_communication_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                                 //              (terminated)
		.av_lock               (),                                                                                                 //              (terminated)
		.av_clken              (),                                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                                             //              (terminated)
		.av_outputenable       ()                                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (15),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) main_memory_communication_s1_translator (
		.clk                   (clk_clk),                                                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                          //                    reset.reset
		.uav_address           (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (main_memory_communication_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (main_memory_communication_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (main_memory_communication_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (main_memory_communication_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (main_memory_communication_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (main_memory_communication_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (main_memory_communication_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                        //              (terminated)
		.av_begintransfer      (),                                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                                        //              (terminated)
		.av_burstcount         (),                                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                                        //              (terminated)
		.av_lock               (),                                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                                    //              (terminated)
		.av_debugaccess        (),                                                                                        //              (terminated)
		.av_outputenable       ()                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_communication_s1_translator (
		.clk                   (clk_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                //                    reset.reset
		.uav_address           (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_communication_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_communication_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_communication_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_communication_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_communication_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_communication_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_communication_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_communication_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_communication_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) descriptor_memory_s1_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (descriptor_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (descriptor_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (descriptor_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (descriptor_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (descriptor_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sgdma_tx_csr_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sgdma_tx_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sgdma_tx_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sgdma_tx_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sgdma_tx_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sgdma_tx_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sgdma_rx_csr_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sgdma_rx_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sgdma_rx_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sgdma_rx_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sgdma_rx_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sgdma_rx_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) tse_mac_control_port_translator (
		.clk                   (clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (tse_mac_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (tse_mac_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (tse_mac_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (tse_mac_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (tse_mac_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_communication_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                       //                    reset.reset
		.uav_address           (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_communication_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                                     //              (terminated)
		.av_byteenable         (),                                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                                     //              (terminated)
		.av_lock               (),                                                                                                     //              (terminated)
		.av_clken              (),                                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                                 //              (terminated)
		.av_debugaccess        (),                                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shared_memory_s1_translator (
		.clk                   (clk_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (shared_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (shared_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (shared_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shared_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (shared_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (shared_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (shared_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mutex_shared_memory_s1_translator (
		.clk                   (clk_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (mutex_shared_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (mutex_shared_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (mutex_shared_memory_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (mutex_shared_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (mutex_shared_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (mutex_shared_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) interval_timer_s1_translator (
		.clk                   (clk_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address           (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (interval_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (interval_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (interval_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (interval_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (interval_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_communication_led_s1_translator (
		.clk                   (clk_clk),                                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address           (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_communication_led_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pio_communication_led_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (pio_communication_led_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pio_communication_led_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (pio_communication_led_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                                    //              (terminated)
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_byteenable         (),                                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shared_memory_s2_translator (
		.clk                   (clk_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (shared_memory_s2_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (shared_memory_s2_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (shared_memory_s2_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shared_memory_s2_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (shared_memory_s2_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (shared_memory_s2_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (shared_memory_s2_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (15),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) main_memory_car_controll_s1_translator (
		.clk                   (clk_clk),                                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address           (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (main_memory_car_controll_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (main_memory_car_controll_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (main_memory_car_controll_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (main_memory_car_controll_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (main_memory_car_controll_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (main_memory_car_controll_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (main_memory_car_controll_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                       //              (terminated)
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_car_controll_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                                         //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                  //                    reset.reset
		.uav_address           (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_car_controll_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                                //              (terminated)
		.av_burstcount         (),                                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                                //              (terminated)
		.av_lock               (),                                                                                                //              (terminated)
		.av_clken              (),                                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                                            //              (terminated)
		.av_outputenable       ()                                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_carcontrol_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                    //                    reset.reset
		.uav_address           (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                                  //              (terminated)
		.av_lock               (),                                                                                                  //              (terminated)
		.av_clken              (),                                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                                   //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) nios2_communication_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                            //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.av_address       (nios2_communication_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_communication_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_communication_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_communication_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_communication_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_communication_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_communication_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_communication_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_communication_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_communication_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_communication_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                                              //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                               //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                                            //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                                      //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                                        //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                               //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) nios2_communication_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                     //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.av_address       (nios2_communication_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_communication_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_communication_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_communication_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_communication_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_communication_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_communication_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_communication_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_communication_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_communication_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_communication_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                                  //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                                   //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                                //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                                          //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                                            //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                                   //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) nios2_car_controll_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                    //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.av_address       (nios2_car_controll_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_car_controll_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_car_controll_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_car_controll_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_car_controll_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_car_controll_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_car_controll_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_car_controll_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_car_controll_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_car_controll_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_car_controll_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_002_src_valid),                                                                 //        rp.valid
		.rp_data          (rsp_xbar_mux_002_src_data),                                                                  //          .data
		.rp_channel       (rsp_xbar_mux_002_src_channel),                                                               //          .channel
		.rp_startofpacket (rsp_xbar_mux_002_src_startofpacket),                                                         //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_002_src_endofpacket),                                                           //          .endofpacket
		.rp_ready         (rsp_xbar_mux_002_src_ready)                                                                  //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                           //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.av_address       (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                                         //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                                          //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                                       //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                                 //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                                   //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                                          //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (4),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_003_src1_valid),                                                        //        rp.valid
		.rp_data          (rsp_xbar_demux_003_src1_data),                                                         //          .data
		.rp_channel       (rsp_xbar_demux_003_src1_channel),                                                      //          .channel
		.rp_startofpacket (rsp_xbar_demux_003_src1_startofpacket),                                                //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),                                                  //          .endofpacket
		.rp_ready         (rsp_xbar_demux_003_src1_ready)                                                         //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (5),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                               //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.av_address       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_003_src2_valid),                                                         //        rp.valid
		.rp_data          (rsp_xbar_demux_003_src2_data),                                                          //          .data
		.rp_channel       (rsp_xbar_demux_003_src2_channel),                                                       //          .channel
		.rp_startofpacket (rsp_xbar_demux_003_src2_startofpacket),                                                 //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_003_src2_endofpacket),                                                   //          .endofpacket
		.rp_ready         (rsp_xbar_demux_003_src2_ready)                                                          //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (6),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                              //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_003_src3_valid),                                                        //        rp.valid
		.rp_data          (rsp_xbar_demux_003_src3_data),                                                         //          .data
		.rp_channel       (rsp_xbar_demux_003_src3_channel),                                                      //          .channel
		.rp_startofpacket (rsp_xbar_demux_003_src3_startofpacket),                                                //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_003_src3_endofpacket),                                                  //          .endofpacket
		.rp_ready         (rsp_xbar_demux_003_src3_ready)                                                         //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (7),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                               //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.av_address       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_003_src4_valid),                                                         //        rp.valid
		.rp_data          (rsp_xbar_demux_003_src4_data),                                                          //          .data
		.rp_channel       (rsp_xbar_demux_003_src4_channel),                                                       //          .channel
		.rp_startofpacket (rsp_xbar_demux_003_src4_startofpacket),                                                 //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_003_src4_endofpacket),                                                   //          .endofpacket
		.rp_ready         (rsp_xbar_demux_003_src4_ready)                                                          //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (8),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_rx_m_write_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                      //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.av_address       (sgdma_rx_m_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_m_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_m_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_m_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_m_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_m_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_001_src2_valid),                                                //        rp.valid
		.rp_data          (rsp_xbar_demux_001_src2_data),                                                 //          .data
		.rp_channel       (rsp_xbar_demux_001_src2_channel),                                              //          .channel
		.rp_startofpacket (rsp_xbar_demux_001_src2_startofpacket),                                        //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),                                          //          .endofpacket
		.rp_ready         (rsp_xbar_demux_001_src2_ready)                                                 //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (9),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_tx_m_read_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                     //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address       (sgdma_tx_m_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_m_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_m_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_m_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_m_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_m_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_001_src3_valid),                                               //        rp.valid
		.rp_data          (rsp_xbar_demux_001_src3_data),                                                //          .data
		.rp_channel       (rsp_xbar_demux_001_src3_channel),                                             //          .channel
		.rp_startofpacket (rsp_xbar_demux_001_src3_startofpacket),                                       //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_001_src3_endofpacket),                                         //          .endofpacket
		.rp_ready         (rsp_xbar_demux_001_src3_ready)                                                //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                             //       clk_reset.reset
		.m0_address              (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                                   //                .channel
		.rf_sink_ready           (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                             // clk_reset.reset
		.in_data           (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) main_memory_communication_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                                        //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                                        //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                         //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                                      //                .channel
		.rf_sink_ready           (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_communication_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_communication_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                                //                .channel
		.rf_sink_ready           (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) descriptor_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                              //                .channel
		.rf_sink_ready           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sgdma_tx_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                   //                .channel
		.rf_sink_ready           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sgdma_rx_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                   //                .channel
		.rf_sink_ready           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) tse_mac_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                           //                .channel
		.rf_sink_ready           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                                                //                .channel
		.rf_sink_ready           (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                 // clk_reset.reset
		.in_data           (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                                           // (terminated)
		.csr_readdata      (),                                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                           // (terminated)
		.almost_full_data  (),                                                                                                               // (terminated)
		.almost_empty_data (),                                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                                           // (terminated)
		.out_empty         (),                                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                                           // (terminated)
		.out_error         (),                                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                                           // (terminated)
		.out_channel       ()                                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shared_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                       //                .channel
		.rf_sink_ready           (shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_009_src_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_009_src_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_009_src_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_009_src_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_009_src_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_009_src_channel),                                                                //                .channel
		.rf_sink_ready           (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) interval_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_010_src_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_010_src_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_010_src_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_010_src_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_010_src_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_010_src_channel),                                                           //                .channel
		.rf_sink_ready           (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_communication_led_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                              //                .channel
		.rf_sink_ready           (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shared_memory_s2_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shared_memory_s2_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src2_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src2_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_002_src2_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src2_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src2_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src2_channel),                                                       //                .channel
		.rf_sink_ready           (shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shared_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shared_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shared_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shared_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shared_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shared_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shared_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shared_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_013_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_013_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_013_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_013_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_013_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_013_src_channel),                                                                     //                .channel
		.rf_sink_ready           (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                            //       clk_reset.reset
		.m0_address              (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_014_src_ready),                                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_014_src_valid),                                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_014_src_data),                                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_014_src_startofpacket),                                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_014_src_endofpacket),                                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_014_src_channel),                                                                              //                .channel
		.rf_sink_ready           (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                            // clk_reset.reset
		.in_data           (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                                      // (terminated)
		.csr_readdata      (),                                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                      // (terminated)
		.almost_full_data  (),                                                                                                          // (terminated)
		.almost_empty_data (),                                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                                      // (terminated)
		.out_empty         (),                                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                                      // (terminated)
		.out_error         (),                                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                                      // (terminated)
		.out_channel       ()                                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                              //       clk_reset.reset
		.m0_address              (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_002_src5_ready),                                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_002_src5_valid),                                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_002_src5_data),                                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_002_src5_startofpacket),                                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_002_src5_endofpacket),                                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_002_src5_channel),                                                                             //                .channel
		.rf_sink_ready           (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                              // clk_reset.reset
		.in_data           (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                                        // (terminated)
		.csr_readdata      (),                                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                        // (terminated)
		.almost_full_data  (),                                                                                                            // (terminated)
		.almost_empty_data (),                                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                                        // (terminated)
		.out_empty         (),                                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                                        // (terminated)
		.out_error         (),                                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                                        // (terminated)
		.out_channel       ()                                                                                                             // (terminated)
	);

	nios_system_addr_router addr_router (
		.sink_ready         (nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_communication_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                                              //          .valid
		.src_data           (addr_router_src_data),                                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                         //          .endofpacket
	);

	nios_system_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_communication_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                              //          .endofpacket
	);

	nios_system_addr_router_002 addr_router_002 (
		.sink_ready         (nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_car_controll_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                                  //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                                  //          .valid
		.src_data           (addr_router_002_src_data),                                                                   //          .data
		.src_channel        (addr_router_002_src_channel),                                                                //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                             //          .endofpacket
	);

	nios_system_addr_router_003 addr_router_003 (
		.sink_ready         (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_car_controll_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                                         //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                                         //          .valid
		.src_data           (addr_router_003_src_data),                                                                          //          .data
		.src_channel        (addr_router_003_src_channel),                                                                       //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                                    //          .endofpacket
	);

	nios_system_addr_router_004 addr_router_004 (
		.sink_ready         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                            //          .valid
		.src_data           (addr_router_004_src_data),                                                             //          .data
		.src_channel        (addr_router_004_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                       //          .endofpacket
	);

	nios_system_addr_router_004 addr_router_005 (
		.sink_ready         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                             //          .valid
		.src_data           (addr_router_005_src_data),                                                              //          .data
		.src_channel        (addr_router_005_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                        //          .endofpacket
	);

	nios_system_addr_router_004 addr_router_006 (
		.sink_ready         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_006_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_006_src_valid),                                                            //          .valid
		.src_data           (addr_router_006_src_data),                                                             //          .data
		.src_channel        (addr_router_006_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_006_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_006_src_endofpacket)                                                       //          .endofpacket
	);

	nios_system_addr_router_004 addr_router_007 (
		.sink_ready         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (addr_router_007_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_007_src_valid),                                                             //          .valid
		.src_data           (addr_router_007_src_data),                                                              //          .data
		.src_channel        (addr_router_007_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_007_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_007_src_endofpacket)                                                        //          .endofpacket
	);

	nios_system_addr_router_008 addr_router_008 (
		.sink_ready         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (addr_router_008_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_008_src_valid),                                                    //          .valid
		.src_data           (addr_router_008_src_data),                                                     //          .data
		.src_channel        (addr_router_008_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_008_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_008_src_endofpacket)                                               //          .endofpacket
	);

	nios_system_addr_router_008 addr_router_009 (
		.sink_ready         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_009_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_009_src_valid),                                                   //          .valid
		.src_data           (addr_router_009_src_data),                                                    //          .data
		.src_channel        (addr_router_009_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_009_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_009_src_endofpacket)                                              //          .endofpacket
	);

	nios_system_id_router id_router (
		.sink_ready         (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_communication_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                                              //          .valid
		.src_data           (id_router_src_data),                                                                               //          .data
		.src_channel        (id_router_src_channel),                                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                         //          .endofpacket
	);

	nios_system_id_router_001 id_router_001 (
		.sink_ready         (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (main_memory_communication_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                                 //       src.ready
		.src_valid          (id_router_001_src_valid),                                                                 //          .valid
		.src_data           (id_router_001_src_data),                                                                  //          .data
		.src_channel        (id_router_001_src_channel),                                                               //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                            //          .endofpacket
	);

	nios_system_id_router id_router_002 (
		.sink_ready         (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_communication_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                           //       src.ready
		.src_valid          (id_router_002_src_valid),                                                           //          .valid
		.src_data           (id_router_002_src_data),                                                            //          .data
		.src_channel        (id_router_002_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                      //          .endofpacket
	);

	nios_system_id_router_003 id_router_003 (
		.sink_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                         //       src.ready
		.src_valid          (id_router_003_src_valid),                                                         //          .valid
		.src_data           (id_router_003_src_data),                                                          //          .data
		.src_channel        (id_router_003_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                    //          .endofpacket
	);

	nios_system_id_router_004 id_router_004 (
		.sink_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                 //       src.ready
		.src_valid          (id_router_004_src_valid),                                                 //          .valid
		.src_data           (id_router_004_src_data),                                                  //          .data
		.src_channel        (id_router_004_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                            //          .endofpacket
	);

	nios_system_id_router_004 id_router_005 (
		.sink_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                 //       src.ready
		.src_valid          (id_router_005_src_valid),                                                 //          .valid
		.src_data           (id_router_005_src_data),                                                  //          .data
		.src_channel        (id_router_005_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                            //          .endofpacket
	);

	nios_system_id_router_004 id_router_006 (
		.sink_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                         //       src.ready
		.src_valid          (id_router_006_src_valid),                                                         //          .valid
		.src_data           (id_router_006_src_data),                                                          //          .data
		.src_channel        (id_router_006_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                    //          .endofpacket
	);

	nios_system_id_router_004 id_router_007 (
		.sink_ready         (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_communication_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                       // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                                              //       src.ready
		.src_valid          (id_router_007_src_valid),                                                                              //          .valid
		.src_data           (id_router_007_src_data),                                                                               //          .data
		.src_channel        (id_router_007_src_channel),                                                                            //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                                      //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                                         //          .endofpacket
	);

	nios_system_id_router_004 id_router_008 (
		.sink_ready         (shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                     //       src.ready
		.src_valid          (id_router_008_src_valid),                                                     //          .valid
		.src_data           (id_router_008_src_data),                                                      //          .data
		.src_channel        (id_router_008_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                //          .endofpacket
	);

	nios_system_id_router_009 id_router_009 (
		.sink_ready         (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mutex_shared_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                           //       src.ready
		.src_valid          (id_router_009_src_valid),                                                           //          .valid
		.src_data           (id_router_009_src_data),                                                            //          .data
		.src_channel        (id_router_009_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                      //          .endofpacket
	);

	nios_system_id_router_009 id_router_010 (
		.sink_ready         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                      //       src.ready
		.src_valid          (id_router_010_src_valid),                                                      //          .valid
		.src_data           (id_router_010_src_data),                                                       //          .data
		.src_channel        (id_router_010_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                 //          .endofpacket
	);

	nios_system_id_router_004 id_router_011 (
		.sink_ready         (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_communication_led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                             //       src.ready
		.src_valid          (id_router_011_src_valid),                                                             //          .valid
		.src_data           (id_router_011_src_data),                                                              //          .data
		.src_channel        (id_router_011_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                        //          .endofpacket
	);

	nios_system_id_router_012 id_router_012 (
		.sink_ready         (shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shared_memory_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                     //       src.ready
		.src_valid          (id_router_012_src_valid),                                                     //          .valid
		.src_data           (id_router_012_src_data),                                                      //          .data
		.src_channel        (id_router_012_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                //          .endofpacket
	);

	nios_system_id_router_013 id_router_013 (
		.sink_ready         (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (main_memory_car_controll_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                                //       src.ready
		.src_valid          (id_router_013_src_valid),                                                                //          .valid
		.src_data           (id_router_013_src_data),                                                                 //          .data
		.src_channel        (id_router_013_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                           //          .endofpacket
	);

	nios_system_id_router_013 id_router_014 (
		.sink_ready         (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_car_controll_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                                         //       src.ready
		.src_valid          (id_router_014_src_valid),                                                                         //          .valid
		.src_data           (id_router_014_src_data),                                                                          //          .data
		.src_channel        (id_router_014_src_channel),                                                                       //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                                    //          .endofpacket
	);

	nios_system_id_router_012 id_router_015 (
		.sink_ready         (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_carcontrol_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                                           //       src.ready
		.src_valid          (id_router_015_src_valid),                                                                           //          .valid
		.src_data           (id_router_015_src_data),                                                                            //          .data
		.src_channel        (id_router_015_src_channel),                                                                         //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                                                   //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                                      //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.VALID_WIDTH               (16),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.VALID_WIDTH               (16),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_003_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_003_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_003_src_data),           //          .data
		.cmd_sink_channel       (addr_router_003_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_003_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_003_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_003_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_003_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_003_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_003_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_003_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_003_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                                    // reset_in0.reset
		.reset_in1  (nios2_communication_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (nios2_car_controll_jtag_debug_module_reset_reset),  // reset_in2.reset
		.clk        (clk_clk),                                           //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),                    // reset_out.reset
		.reset_in3  (1'b0),                                              // (terminated)
		.reset_in4  (1'b0),                                              // (terminated)
		.reset_in5  (1'b0),                                              // (terminated)
		.reset_in6  (1'b0),                                              // (terminated)
		.reset_in7  (1'b0),                                              // (terminated)
		.reset_in8  (1'b0),                                              // (terminated)
		.reset_in9  (1'b0),                                              // (terminated)
		.reset_in10 (1'b0),                                              // (terminated)
		.reset_in11 (1'b0),                                              // (terminated)
		.reset_in12 (1'b0),                                              // (terminated)
		.reset_in13 (1'b0),                                              // (terminated)
		.reset_in14 (1'b0),                                              // (terminated)
		.reset_in15 (1'b0)                                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //           .endofpacket
	);

	nios_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_002_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_002_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_002_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_002_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_002_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_002_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_002_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_002_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_002_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_002_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_002_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_002_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_002_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_002_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_002_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_002_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_002_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_002_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_002_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_002_src5_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_003_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_003_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_003_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_003_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket)    //           .endofpacket
	);

	nios_system_cmd_xbar_demux_004 cmd_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 cmd_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_005_src_ready),             //      sink.ready
		.sink_channel       (addr_router_005_src_channel),           //          .channel
		.sink_data          (addr_router_005_src_data),              //          .data
		.sink_startofpacket (addr_router_005_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_005_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_005_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 cmd_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_006_src_ready),             //      sink.ready
		.sink_channel       (addr_router_006_src_channel),           //          .channel
		.sink_data          (addr_router_006_src_data),              //          .data
		.sink_startofpacket (addr_router_006_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_006_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_006_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 cmd_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_007_src_ready),             //      sink.ready
		.sink_channel       (addr_router_007_src_channel),           //          .channel
		.sink_data          (addr_router_007_src_data),              //          .data
		.sink_startofpacket (addr_router_007_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_007_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_007_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 cmd_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_008_src_ready),             //      sink.ready
		.sink_channel       (addr_router_008_src_channel),           //          .channel
		.sink_data          (addr_router_008_src_data),              //          .data
		.sink_startofpacket (addr_router_008_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_008_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_008_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 cmd_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_009_src_ready),             //      sink.ready
		.sink_channel       (addr_router_009_src_channel),           //          .channel
		.sink_data          (addr_router_009_src_data),              //          .data
		.sink_startofpacket (addr_router_009_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_009_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_009_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_008_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_008_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_008_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_008_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_009_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_009_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_009_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_009_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_003 cmd_xbar_mux_003 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src3_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_004_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_005_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_006_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_006_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_006_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_006_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (cmd_xbar_demux_007_src0_ready),         //     sink4.ready
		.sink4_valid         (cmd_xbar_demux_007_src0_valid),         //          .valid
		.sink4_channel       (cmd_xbar_demux_007_src0_channel),       //          .channel
		.sink4_data          (cmd_xbar_demux_007_src0_data),          //          .data
		.sink4_startofpacket (cmd_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (cmd_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_009 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_009_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_009_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_009_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src9_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src9_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src9_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src9_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src9_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src9_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_010 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_010_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_010_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_010_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_010_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_010_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_010_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src10_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src1_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src1_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src1_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_002_src1_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src1_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket)     //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_013 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_013_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_013_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_013_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_013_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_013_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_013_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src3_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src3_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src3_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src3_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_014 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_014_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_014_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_014_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_014_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_014_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_014_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src4_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src4_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src4_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src4_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src4_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src4_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_003_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_003_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_003_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_003_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_003_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_003_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_003_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_003_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_003_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_003_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_003_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_003_src3_endofpacket),   //          .endofpacket
		.src4_ready         (rsp_xbar_demux_003_src4_ready),         //      src4.ready
		.src4_valid         (rsp_xbar_demux_003_src4_valid),         //          .valid
		.src4_data          (rsp_xbar_demux_003_src4_data),          //          .data
		.src4_channel       (rsp_xbar_demux_003_src4_channel),       //          .channel
		.src4_startofpacket (rsp_xbar_demux_003_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (rsp_xbar_demux_003_src4_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_009_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_010_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_013 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_013_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_013_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_014 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_014_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_014_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_014_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_014_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_014_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_014_src1_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_004 rsp_xbar_demux_015 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_009_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_010_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_012_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_013_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_014_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_015_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux_003 rsp_xbar_mux_003 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_013_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_013_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_014_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_014_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_014_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_014_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_014_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_014_src1_endofpacket)    //          .endofpacket
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_communication_d_irq_irq)   //    sender.irq
	);

	nios_system_irq_mapper_001 irq_mapper_001 (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),   // receiver0.irq
		.sender_irq    (nios2_car_controll_d_irq_irq)    //    sender.irq
	);

endmodule
