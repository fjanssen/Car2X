// ethernet_system.v

// Generated using ACDS version 12.1 177 at 2014.06.30.20:20:02

`timescale 1 ps / 1 ps
module ethernet_system (
		input  wire        ethernet_subsys_clk_in_clk,        //   ethernet_subsys_clk_in.clk
		output wire        ethernet_bridge_s0_waitrequest,    //       ethernet_bridge_s0.waitrequest
		output wire [31:0] ethernet_bridge_s0_readdata,       //                         .readdata
		output wire        ethernet_bridge_s0_readdatavalid,  //                         .readdatavalid
		input  wire [0:0]  ethernet_bridge_s0_burstcount,     //                         .burstcount
		input  wire [31:0] ethernet_bridge_s0_writedata,      //                         .writedata
		input  wire [10:0] ethernet_bridge_s0_address,        //                         .address
		input  wire        ethernet_bridge_s0_write,          //                         .write
		input  wire        ethernet_bridge_s0_read,           //                         .read
		input  wire [3:0]  ethernet_bridge_s0_byteenable,     //                         .byteenable
		input  wire        ethernet_bridge_s0_debugaccess,    //                         .debugaccess
		input  wire        sgdma_rx_m_write_waitrequest,      //         sgdma_rx_m_write.waitrequest
		output wire [31:0] sgdma_rx_m_write_address,          //                         .address
		output wire        sgdma_rx_m_write_write,            //                         .write
		output wire [31:0] sgdma_rx_m_write_writedata,        //                         .writedata
		output wire [3:0]  sgdma_rx_m_write_byteenable,       //                         .byteenable
		input  wire [3:0]  tse_conduit_connection_rgmii_in,   //   tse_conduit_connection.rgmii_in
		output wire [3:0]  tse_conduit_connection_rgmii_out,  //                         .rgmii_out
		input  wire        tse_conduit_connection_rx_control, //                         .rx_control
		output wire        tse_conduit_connection_tx_control, //                         .tx_control
		input  wire        tse_conduit_connection_tx_clk,     //                         .tx_clk
		input  wire        tse_conduit_connection_rx_clk,     //                         .rx_clk
		input  wire        tse_conduit_connection_set_10,     //                         .set_10
		input  wire        tse_conduit_connection_set_1000,   //                         .set_1000
		output wire        tse_conduit_connection_ena_10,     //                         .ena_10
		output wire        tse_conduit_connection_eth_mode,   //                         .eth_mode
		output wire        tse_conduit_connection_mdio_out,   //                         .mdio_out
		output wire        tse_conduit_connection_mdio_oen,   //                         .mdio_oen
		input  wire        tse_conduit_connection_mdio_in,    //                         .mdio_in
		output wire        tse_conduit_connection_mdc,        //                         .mdc
		output wire        sgdma_rx_csr_irq_irq,              //         sgdma_rx_csr_irq.irq
		input  wire [31:0] sgdma_tx_m_read_readdata,          //          sgdma_tx_m_read.readdata
		input  wire        sgdma_tx_m_read_readdatavalid,     //                         .readdatavalid
		input  wire        sgdma_tx_m_read_waitrequest,       //                         .waitrequest
		output wire [31:0] sgdma_tx_m_read_address,           //                         .address
		output wire        sgdma_tx_m_read_read,              //                         .read
		output wire        sgdma_tx_csr_irq_irq,              //         sgdma_tx_csr_irq.irq
		input  wire [10:0] descriptor_memory_s2_address,      //     descriptor_memory_s2.address
		input  wire        descriptor_memory_s2_chipselect,   //                         .chipselect
		input  wire        descriptor_memory_s2_clken,        //                         .clken
		output wire [31:0] descriptor_memory_s2_readdata,     //                         .readdata
		input  wire        descriptor_memory_s2_write,        //                         .write
		input  wire [31:0] descriptor_memory_s2_writedata,    //                         .writedata
		input  wire [3:0]  descriptor_memory_s2_byteenable,   //                         .byteenable
		input  wire        ethernet_subsys_reset_in_reset_n   // ethernet_subsys_reset_in.reset_n
	);

	wire          tse_mac_receive_endofpacket;                                                               // tse_mac:ff_rx_eop -> sgdma_rx:in_endofpacket
	wire          tse_mac_receive_valid;                                                                     // tse_mac:ff_rx_dval -> sgdma_rx:in_valid
	wire          tse_mac_receive_startofpacket;                                                             // tse_mac:ff_rx_sop -> sgdma_rx:in_startofpacket
	wire    [5:0] tse_mac_receive_error;                                                                     // tse_mac:rx_err -> sgdma_rx:in_error
	wire    [1:0] tse_mac_receive_empty;                                                                     // tse_mac:ff_rx_mod -> sgdma_rx:in_empty
	wire   [31:0] tse_mac_receive_data;                                                                      // tse_mac:ff_rx_data -> sgdma_rx:in_data
	wire          tse_mac_receive_ready;                                                                     // sgdma_rx:in_ready -> tse_mac:ff_rx_rdy
	wire          sgdma_tx_out_endofpacket;                                                                  // sgdma_tx:out_endofpacket -> tse_mac:ff_tx_eop
	wire          sgdma_tx_out_valid;                                                                        // sgdma_tx:out_valid -> tse_mac:ff_tx_wren
	wire          sgdma_tx_out_startofpacket;                                                                // sgdma_tx:out_startofpacket -> tse_mac:ff_tx_sop
	wire          sgdma_tx_out_error;                                                                        // sgdma_tx:out_error -> tse_mac:ff_tx_err
	wire    [1:0] sgdma_tx_out_empty;                                                                        // sgdma_tx:out_empty -> tse_mac:ff_tx_mod
	wire   [31:0] sgdma_tx_out_data;                                                                         // sgdma_tx:out_data -> tse_mac:ff_tx_data
	wire          sgdma_tx_out_ready;                                                                        // tse_mac:ff_tx_rdy -> sgdma_tx:out_ready
	wire    [0:0] ethernet_bridge_m0_burstcount;                                                             // ethernet_bridge:m0_burstcount -> ethernet_bridge_m0_translator:av_burstcount
	wire          ethernet_bridge_m0_waitrequest;                                                            // ethernet_bridge_m0_translator:av_waitrequest -> ethernet_bridge:m0_waitrequest
	wire   [10:0] ethernet_bridge_m0_address;                                                                // ethernet_bridge:m0_address -> ethernet_bridge_m0_translator:av_address
	wire   [31:0] ethernet_bridge_m0_writedata;                                                              // ethernet_bridge:m0_writedata -> ethernet_bridge_m0_translator:av_writedata
	wire          ethernet_bridge_m0_write;                                                                  // ethernet_bridge:m0_write -> ethernet_bridge_m0_translator:av_write
	wire          ethernet_bridge_m0_read;                                                                   // ethernet_bridge:m0_read -> ethernet_bridge_m0_translator:av_read
	wire   [31:0] ethernet_bridge_m0_readdata;                                                               // ethernet_bridge_m0_translator:av_readdata -> ethernet_bridge:m0_readdata
	wire          ethernet_bridge_m0_debugaccess;                                                            // ethernet_bridge:m0_debugaccess -> ethernet_bridge_m0_translator:av_debugaccess
	wire    [3:0] ethernet_bridge_m0_byteenable;                                                             // ethernet_bridge:m0_byteenable -> ethernet_bridge_m0_translator:av_byteenable
	wire          ethernet_bridge_m0_readdatavalid;                                                          // ethernet_bridge_m0_translator:av_readdatavalid -> ethernet_bridge:m0_readdatavalid
	wire          tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest;                           // tse_mac:waitrequest -> tse_mac_control_port_translator:av_waitrequest
	wire   [31:0] tse_mac_control_port_translator_avalon_anti_slave_0_writedata;                             // tse_mac_control_port_translator:av_writedata -> tse_mac:writedata
	wire    [7:0] tse_mac_control_port_translator_avalon_anti_slave_0_address;                               // tse_mac_control_port_translator:av_address -> tse_mac:address
	wire          tse_mac_control_port_translator_avalon_anti_slave_0_write;                                 // tse_mac_control_port_translator:av_write -> tse_mac:write
	wire          tse_mac_control_port_translator_avalon_anti_slave_0_read;                                  // tse_mac_control_port_translator:av_read -> tse_mac:read
	wire   [31:0] tse_mac_control_port_translator_avalon_anti_slave_0_readdata;                              // tse_mac:readdata -> tse_mac_control_port_translator:av_readdata
	wire   [31:0] sgdma_rx_csr_translator_avalon_anti_slave_0_writedata;                                     // sgdma_rx_csr_translator:av_writedata -> sgdma_rx:csr_writedata
	wire    [3:0] sgdma_rx_csr_translator_avalon_anti_slave_0_address;                                       // sgdma_rx_csr_translator:av_address -> sgdma_rx:csr_address
	wire          sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect;                                    // sgdma_rx_csr_translator:av_chipselect -> sgdma_rx:csr_chipselect
	wire          sgdma_rx_csr_translator_avalon_anti_slave_0_write;                                         // sgdma_rx_csr_translator:av_write -> sgdma_rx:csr_write
	wire          sgdma_rx_csr_translator_avalon_anti_slave_0_read;                                          // sgdma_rx_csr_translator:av_read -> sgdma_rx:csr_read
	wire   [31:0] sgdma_rx_csr_translator_avalon_anti_slave_0_readdata;                                      // sgdma_rx:csr_readdata -> sgdma_rx_csr_translator:av_readdata
	wire   [31:0] sgdma_tx_csr_translator_avalon_anti_slave_0_writedata;                                     // sgdma_tx_csr_translator:av_writedata -> sgdma_tx:csr_writedata
	wire    [3:0] sgdma_tx_csr_translator_avalon_anti_slave_0_address;                                       // sgdma_tx_csr_translator:av_address -> sgdma_tx:csr_address
	wire          sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect;                                    // sgdma_tx_csr_translator:av_chipselect -> sgdma_tx:csr_chipselect
	wire          sgdma_tx_csr_translator_avalon_anti_slave_0_write;                                         // sgdma_tx_csr_translator:av_write -> sgdma_tx:csr_write
	wire          sgdma_tx_csr_translator_avalon_anti_slave_0_read;                                          // sgdma_tx_csr_translator:av_read -> sgdma_tx:csr_read
	wire   [31:0] sgdma_tx_csr_translator_avalon_anti_slave_0_readdata;                                      // sgdma_tx:csr_readdata -> sgdma_tx_csr_translator:av_readdata
	wire          sgdma_rx_descriptor_read_waitrequest;                                                      // sgdma_rx_descriptor_read_translator:av_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	wire   [31:0] sgdma_rx_descriptor_read_address;                                                          // sgdma_rx:descriptor_read_address -> sgdma_rx_descriptor_read_translator:av_address
	wire          sgdma_rx_descriptor_read_read;                                                             // sgdma_rx:descriptor_read_read -> sgdma_rx_descriptor_read_translator:av_read
	wire   [31:0] sgdma_rx_descriptor_read_readdata;                                                         // sgdma_rx_descriptor_read_translator:av_readdata -> sgdma_rx:descriptor_read_readdata
	wire          sgdma_rx_descriptor_read_readdatavalid;                                                    // sgdma_rx_descriptor_read_translator:av_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	wire          sgdma_rx_descriptor_write_waitrequest;                                                     // sgdma_rx_descriptor_write_translator:av_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	wire   [31:0] sgdma_rx_descriptor_write_writedata;                                                       // sgdma_rx:descriptor_write_writedata -> sgdma_rx_descriptor_write_translator:av_writedata
	wire   [31:0] sgdma_rx_descriptor_write_address;                                                         // sgdma_rx:descriptor_write_address -> sgdma_rx_descriptor_write_translator:av_address
	wire          sgdma_rx_descriptor_write_write;                                                           // sgdma_rx:descriptor_write_write -> sgdma_rx_descriptor_write_translator:av_write
	wire          sgdma_tx_descriptor_read_waitrequest;                                                      // sgdma_tx_descriptor_read_translator:av_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	wire   [31:0] sgdma_tx_descriptor_read_address;                                                          // sgdma_tx:descriptor_read_address -> sgdma_tx_descriptor_read_translator:av_address
	wire          sgdma_tx_descriptor_read_read;                                                             // sgdma_tx:descriptor_read_read -> sgdma_tx_descriptor_read_translator:av_read
	wire   [31:0] sgdma_tx_descriptor_read_readdata;                                                         // sgdma_tx_descriptor_read_translator:av_readdata -> sgdma_tx:descriptor_read_readdata
	wire          sgdma_tx_descriptor_read_readdatavalid;                                                    // sgdma_tx_descriptor_read_translator:av_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	wire          sgdma_tx_descriptor_write_waitrequest;                                                     // sgdma_tx_descriptor_write_translator:av_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	wire   [31:0] sgdma_tx_descriptor_write_writedata;                                                       // sgdma_tx:descriptor_write_writedata -> sgdma_tx_descriptor_write_translator:av_writedata
	wire   [31:0] sgdma_tx_descriptor_write_address;                                                         // sgdma_tx:descriptor_write_address -> sgdma_tx_descriptor_write_translator:av_address
	wire          sgdma_tx_descriptor_write_write;                                                           // sgdma_tx:descriptor_write_write -> sgdma_tx_descriptor_write_translator:av_write
	wire   [31:0] descriptor_memory_s1_translator_avalon_anti_slave_0_writedata;                             // descriptor_memory_s1_translator:av_writedata -> descriptor_memory:writedata
	wire   [10:0] descriptor_memory_s1_translator_avalon_anti_slave_0_address;                               // descriptor_memory_s1_translator:av_address -> descriptor_memory:address
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect;                            // descriptor_memory_s1_translator:av_chipselect -> descriptor_memory:chipselect
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_clken;                                 // descriptor_memory_s1_translator:av_clken -> descriptor_memory:clken
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_write;                                 // descriptor_memory_s1_translator:av_write -> descriptor_memory:write
	wire   [31:0] descriptor_memory_s1_translator_avalon_anti_slave_0_readdata;                              // descriptor_memory:readdata -> descriptor_memory_s1_translator:av_readdata
	wire    [3:0] descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable;                            // descriptor_memory_s1_translator:av_byteenable -> descriptor_memory:byteenable
	wire          ethernet_bridge_m0_translator_avalon_universal_master_0_waitrequest;                       // ethernet_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> ethernet_bridge_m0_translator:uav_waitrequest
	wire    [2:0] ethernet_bridge_m0_translator_avalon_universal_master_0_burstcount;                        // ethernet_bridge_m0_translator:uav_burstcount -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] ethernet_bridge_m0_translator_avalon_universal_master_0_writedata;                         // ethernet_bridge_m0_translator:uav_writedata -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [10:0] ethernet_bridge_m0_translator_avalon_universal_master_0_address;                           // ethernet_bridge_m0_translator:uav_address -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          ethernet_bridge_m0_translator_avalon_universal_master_0_lock;                              // ethernet_bridge_m0_translator:uav_lock -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          ethernet_bridge_m0_translator_avalon_universal_master_0_write;                             // ethernet_bridge_m0_translator:uav_write -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          ethernet_bridge_m0_translator_avalon_universal_master_0_read;                              // ethernet_bridge_m0_translator:uav_read -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] ethernet_bridge_m0_translator_avalon_universal_master_0_readdata;                          // ethernet_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> ethernet_bridge_m0_translator:uav_readdata
	wire          ethernet_bridge_m0_translator_avalon_universal_master_0_debugaccess;                       // ethernet_bridge_m0_translator:uav_debugaccess -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] ethernet_bridge_m0_translator_avalon_universal_master_0_byteenable;                        // ethernet_bridge_m0_translator:uav_byteenable -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          ethernet_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                     // ethernet_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> ethernet_bridge_m0_translator:uav_readdatavalid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // tse_mac_control_port_translator:uav_waitrequest -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;              // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> tse_mac_control_port_translator:uav_burstcount
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;               // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> tse_mac_control_port_translator:uav_writedata
	wire   [10:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address;                 // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_address -> tse_mac_control_port_translator:uav_address
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write;                   // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_write -> tse_mac_control_port_translator:uav_write
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                    // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> tse_mac_control_port_translator:uav_lock
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read;                    // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_read -> tse_mac_control_port_translator:uav_read
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                // tse_mac_control_port_translator:uav_readdata -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // tse_mac_control_port_translator:uav_readdatavalid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> tse_mac_control_port_translator:uav_debugaccess
	wire    [3:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;              // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> tse_mac_control_port_translator:uav_byteenable
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;            // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;             // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;            // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // sgdma_rx_csr_translator:uav_waitrequest -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_rx_csr_translator:uav_burstcount
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                       // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_rx_csr_translator:uav_writedata
	wire   [10:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address;                         // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_rx_csr_translator:uav_address
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write;                           // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_rx_csr_translator:uav_write
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock;                            // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_rx_csr_translator:uav_lock
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read;                            // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_rx_csr_translator:uav_read
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                        // sgdma_rx_csr_translator:uav_readdata -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // sgdma_rx_csr_translator:uav_readdatavalid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_rx_csr_translator:uav_debugaccess
	wire    [3:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_rx_csr_translator:uav_byteenable
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                     // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // sgdma_tx_csr_translator:uav_waitrequest -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_tx_csr_translator:uav_burstcount
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                       // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_tx_csr_translator:uav_writedata
	wire   [10:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address;                         // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_tx_csr_translator:uav_address
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write;                           // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_tx_csr_translator:uav_write
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock;                            // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_tx_csr_translator:uav_lock
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read;                            // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_tx_csr_translator:uav_read
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                        // sgdma_tx_csr_translator:uav_readdata -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // sgdma_tx_csr_translator:uav_readdatavalid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_tx_csr_translator:uav_debugaccess
	wire    [3:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_tx_csr_translator:uav_byteenable
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                     // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest;                 // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_descriptor_read_translator:uav_waitrequest
	wire    [2:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount;                  // sgdma_rx_descriptor_read_translator:uav_burstcount -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata;                   // sgdma_rx_descriptor_read_translator:uav_writedata -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address;                     // sgdma_rx_descriptor_read_translator:uav_address -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock;                        // sgdma_rx_descriptor_read_translator:uav_lock -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write;                       // sgdma_rx_descriptor_read_translator:uav_write -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read;                        // sgdma_rx_descriptor_read_translator:uav_read -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata;                    // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_descriptor_read_translator:uav_readdata
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess;                 // sgdma_rx_descriptor_read_translator:uav_debugaccess -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable;                  // sgdma_rx_descriptor_read_translator:uav_byteenable -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid;               // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_descriptor_read_translator:uav_readdatavalid
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest;                // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_descriptor_write_translator:uav_waitrequest
	wire    [2:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount;                 // sgdma_rx_descriptor_write_translator:uav_burstcount -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata;                  // sgdma_rx_descriptor_write_translator:uav_writedata -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address;                    // sgdma_rx_descriptor_write_translator:uav_address -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock;                       // sgdma_rx_descriptor_write_translator:uav_lock -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write;                      // sgdma_rx_descriptor_write_translator:uav_write -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read;                       // sgdma_rx_descriptor_write_translator:uav_read -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata;                   // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_descriptor_write_translator:uav_readdata
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess;                // sgdma_rx_descriptor_write_translator:uav_debugaccess -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable;                 // sgdma_rx_descriptor_write_translator:uav_byteenable -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid;              // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_descriptor_write_translator:uav_readdatavalid
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest;                 // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_descriptor_read_translator:uav_waitrequest
	wire    [2:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount;                  // sgdma_tx_descriptor_read_translator:uav_burstcount -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata;                   // sgdma_tx_descriptor_read_translator:uav_writedata -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address;                     // sgdma_tx_descriptor_read_translator:uav_address -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock;                        // sgdma_tx_descriptor_read_translator:uav_lock -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write;                       // sgdma_tx_descriptor_read_translator:uav_write -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read;                        // sgdma_tx_descriptor_read_translator:uav_read -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata;                    // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_descriptor_read_translator:uav_readdata
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess;                 // sgdma_tx_descriptor_read_translator:uav_debugaccess -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable;                  // sgdma_tx_descriptor_read_translator:uav_byteenable -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid;               // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_descriptor_read_translator:uav_readdatavalid
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest;                // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_descriptor_write_translator:uav_waitrequest
	wire    [2:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount;                 // sgdma_tx_descriptor_write_translator:uav_burstcount -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata;                  // sgdma_tx_descriptor_write_translator:uav_writedata -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address;                    // sgdma_tx_descriptor_write_translator:uav_address -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock;                       // sgdma_tx_descriptor_write_translator:uav_lock -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write;                      // sgdma_tx_descriptor_write_translator:uav_write -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read;                       // sgdma_tx_descriptor_write_translator:uav_read -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata;                   // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_descriptor_write_translator:uav_readdata
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess;                // sgdma_tx_descriptor_write_translator:uav_debugaccess -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable;                 // sgdma_tx_descriptor_write_translator:uav_byteenable -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid;              // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_descriptor_write_translator:uav_readdatavalid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // descriptor_memory_s1_translator:uav_waitrequest -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;              // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> descriptor_memory_s1_translator:uav_burstcount
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;               // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> descriptor_memory_s1_translator:uav_writedata
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                 // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> descriptor_memory_s1_translator:uav_address
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                   // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> descriptor_memory_s1_translator:uav_write
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> descriptor_memory_s1_translator:uav_lock
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> descriptor_memory_s1_translator:uav_read
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                // descriptor_memory_s1_translator:uav_readdata -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // descriptor_memory_s1_translator:uav_readdatavalid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> descriptor_memory_s1_translator:uav_debugaccess
	wire    [3:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;              // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> descriptor_memory_s1_translator:uav_byteenable
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;            // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;             // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;            // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;              // ethernet_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                    // ethernet_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;            // ethernet_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire   [81:0] ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                     // ethernet_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                    // addr_router:sink_ready -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                   // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire   [81:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data;                    // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid;                           // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [81:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data;                            // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_001:sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid;                           // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [81:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data;                            // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_002:sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;        // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;              // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;      // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [102:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;               // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;              // addr_router_001:sink_ready -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;       // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;             // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;     // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [102:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;              // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;             // addr_router_002:sink_ready -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;        // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;              // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;      // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [102:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;               // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;              // addr_router_003:sink_ready -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;       // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;             // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;     // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [102:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;              // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;             // addr_router_004:sink_ready -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                   // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [102:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_003:sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                               // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                     // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                             // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire   [81:0] addr_router_src_data;                                                                      // addr_router:src_data -> limiter:cmd_sink_data
	wire    [2:0] addr_router_src_channel;                                                                   // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                     // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                               // limiter:rsp_src_endofpacket -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                     // limiter:rsp_src_valid -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                             // limiter:rsp_src_startofpacket -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [81:0] limiter_rsp_src_data;                                                                      // limiter:rsp_src_data -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [2:0] limiter_rsp_src_channel;                                                                   // limiter:rsp_src_channel -> ethernet_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                     // ethernet_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          rst_controller_reset_out_reset;                                                            // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_mux_003:reset, descriptor_memory:reset, descriptor_memory:reset2, descriptor_memory_s1_translator:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ethernet_bridge:reset, ethernet_bridge_m0_translator:reset, ethernet_bridge_m0_translator_avalon_universal_master_0_agent:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, limiter:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_mux:reset, sgdma_rx:system_reset_n, sgdma_rx_csr_translator:reset, sgdma_rx_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_rx_descriptor_read_translator:reset, sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_rx_descriptor_write_translator:reset, sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_tx:system_reset_n, sgdma_tx_csr_translator:reset, sgdma_tx_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_tx_descriptor_read_translator:reset, sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_tx_descriptor_write_translator:reset, sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:reset, tse_mac:reset, tse_mac_control_port_translator:reset, tse_mac_control_port_translator_avalon_universal_slave_0_agent:reset, tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                           // cmd_xbar_demux:src0_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                 // cmd_xbar_demux:src0_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                         // cmd_xbar_demux:src0_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] cmd_xbar_demux_src0_data;                                                                  // cmd_xbar_demux:src0_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] cmd_xbar_demux_src0_channel;                                                               // cmd_xbar_demux:src0_channel -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src1_endofpacket;                                                           // cmd_xbar_demux:src1_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                 // cmd_xbar_demux:src1_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                         // cmd_xbar_demux:src1_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] cmd_xbar_demux_src1_data;                                                                  // cmd_xbar_demux:src1_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] cmd_xbar_demux_src1_channel;                                                               // cmd_xbar_demux:src1_channel -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src2_endofpacket;                                                           // cmd_xbar_demux:src2_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                 // cmd_xbar_demux:src2_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                         // cmd_xbar_demux:src2_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] cmd_xbar_demux_src2_data;                                                                  // cmd_xbar_demux:src2_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] cmd_xbar_demux_src2_channel;                                                               // cmd_xbar_demux:src2_channel -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                           // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                 // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                         // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire   [81:0] rsp_xbar_demux_src0_data;                                                                  // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [2:0] rsp_xbar_demux_src0_channel;                                                               // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                 // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                       // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                             // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                     // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire   [81:0] rsp_xbar_demux_001_src0_data;                                                              // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [2:0] rsp_xbar_demux_001_src0_channel;                                                           // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                             // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                       // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                             // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                     // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire   [81:0] rsp_xbar_demux_002_src0_data;                                                              // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire    [2:0] rsp_xbar_demux_002_src0_channel;                                                           // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                             // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                               // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                             // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire   [81:0] limiter_cmd_src_data;                                                                      // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire    [2:0] limiter_cmd_src_channel;                                                                   // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                     // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                              // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                    // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                            // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire   [81:0] rsp_xbar_mux_src_data;                                                                     // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire    [2:0] rsp_xbar_mux_src_channel;                                                                  // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                    // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          cmd_xbar_demux_src0_ready;                                                                 // tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire          id_router_src_endofpacket;                                                                 // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                       // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                               // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire   [81:0] id_router_src_data;                                                                        // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [2:0] id_router_src_channel;                                                                     // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                       // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_demux_src1_ready;                                                                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire          id_router_001_src_endofpacket;                                                             // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                   // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                           // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire   [81:0] id_router_001_src_data;                                                                    // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [2:0] id_router_001_src_channel;                                                                 // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                   // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_src2_ready;                                                                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	wire          id_router_002_src_endofpacket;                                                             // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                   // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                           // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire   [81:0] id_router_002_src_data;                                                                    // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [2:0] id_router_002_src_channel;                                                                 // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                   // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                       // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                             // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                     // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src0_data;                                                              // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux_003:sink0_data
	wire    [3:0] cmd_xbar_demux_001_src0_channel;                                                           // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                             // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                       // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                             // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                     // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [102:0] cmd_xbar_demux_002_src0_data;                                                              // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_003:sink1_data
	wire    [3:0] cmd_xbar_demux_002_src0_channel;                                                           // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                             // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                       // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_003:sink2_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                             // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_003:sink2_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                     // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_003:sink2_startofpacket
	wire  [102:0] cmd_xbar_demux_003_src0_data;                                                              // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_003:sink2_data
	wire    [3:0] cmd_xbar_demux_003_src0_channel;                                                           // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_003:sink2_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                             // cmd_xbar_mux_003:sink2_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                       // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_003:sink3_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                             // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_003:sink3_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                     // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_003:sink3_startofpacket
	wire  [102:0] cmd_xbar_demux_004_src0_data;                                                              // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_003:sink3_data
	wire    [3:0] cmd_xbar_demux_004_src0_channel;                                                           // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_003:sink3_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                             // cmd_xbar_mux_003:sink3_ready -> cmd_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                       // rsp_xbar_demux_003:src0_endofpacket -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                             // rsp_xbar_demux_003:src0_valid -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                     // rsp_xbar_demux_003:src0_startofpacket -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_demux_003_src0_data;                                                              // rsp_xbar_demux_003:src0_data -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] rsp_xbar_demux_003_src0_channel;                                                           // rsp_xbar_demux_003:src0_channel -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                       // rsp_xbar_demux_003:src1_endofpacket -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                             // rsp_xbar_demux_003:src1_valid -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                     // rsp_xbar_demux_003:src1_startofpacket -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_demux_003_src1_data;                                                              // rsp_xbar_demux_003:src1_data -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] rsp_xbar_demux_003_src1_channel;                                                           // rsp_xbar_demux_003:src1_channel -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_003_src2_endofpacket;                                                       // rsp_xbar_demux_003:src2_endofpacket -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_003_src2_valid;                                                             // rsp_xbar_demux_003:src2_valid -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_003_src2_startofpacket;                                                     // rsp_xbar_demux_003:src2_startofpacket -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_demux_003_src2_data;                                                              // rsp_xbar_demux_003:src2_data -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] rsp_xbar_demux_003_src2_channel;                                                           // rsp_xbar_demux_003:src2_channel -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_003_src3_endofpacket;                                                       // rsp_xbar_demux_003:src3_endofpacket -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_003_src3_valid;                                                             // rsp_xbar_demux_003:src3_valid -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_003_src3_startofpacket;                                                     // rsp_xbar_demux_003:src3_startofpacket -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_demux_003_src3_data;                                                              // rsp_xbar_demux_003:src3_data -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] rsp_xbar_demux_003_src3_channel;                                                           // rsp_xbar_demux_003:src3_channel -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          addr_router_001_src_endofpacket;                                                           // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                 // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                         // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [102:0] addr_router_001_src_data;                                                                  // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [3:0] addr_router_001_src_channel;                                                               // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                 // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_demux_003_src0_ready;                                                             // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_003:src0_ready
	wire          addr_router_002_src_endofpacket;                                                           // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                 // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                         // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [102:0] addr_router_002_src_data;                                                                  // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire    [3:0] addr_router_002_src_channel;                                                               // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                 // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_003_src1_ready;                                                             // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_003:src1_ready
	wire          addr_router_003_src_endofpacket;                                                           // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                 // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                         // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [102:0] addr_router_003_src_data;                                                                  // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire    [3:0] addr_router_003_src_channel;                                                               // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                 // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          rsp_xbar_demux_003_src2_ready;                                                             // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_003:src2_ready
	wire          addr_router_004_src_endofpacket;                                                           // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          addr_router_004_src_valid;                                                                 // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire          addr_router_004_src_startofpacket;                                                         // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [102:0] addr_router_004_src_data;                                                                  // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire    [3:0] addr_router_004_src_channel;                                                               // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire          addr_router_004_src_ready;                                                                 // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire          rsp_xbar_demux_003_src3_ready;                                                             // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_003:src3_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                          // cmd_xbar_mux_003:src_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                // cmd_xbar_mux_003:src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                        // cmd_xbar_mux_003:src_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_mux_003_src_data;                                                                 // cmd_xbar_mux_003:src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [3:0] cmd_xbar_mux_003_src_channel;                                                              // cmd_xbar_mux_003:src_channel -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                             // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                   // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                           // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [102:0] id_router_003_src_data;                                                                    // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [3:0] id_router_003_src_channel;                                                                 // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                   // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire    [2:0] limiter_cmd_valid_data;                                                                    // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (11),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) ethernet_bridge (
		.clk              (ethernet_subsys_clk_in_clk),       //   clk.clk
		.reset            (rst_controller_reset_out_reset),   // reset.reset
		.s0_waitrequest   (ethernet_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (ethernet_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (ethernet_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (ethernet_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (ethernet_bridge_s0_writedata),     //      .writedata
		.s0_address       (ethernet_bridge_s0_address),       //      .address
		.s0_write         (ethernet_bridge_s0_write),         //      .write
		.s0_read          (ethernet_bridge_s0_read),          //      .read
		.s0_byteenable    (ethernet_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (ethernet_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (ethernet_bridge_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (ethernet_bridge_m0_readdata),      //      .readdata
		.m0_readdatavalid (ethernet_bridge_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (ethernet_bridge_m0_burstcount),    //      .burstcount
		.m0_writedata     (ethernet_bridge_m0_writedata),     //      .writedata
		.m0_address       (ethernet_bridge_m0_address),       //      .address
		.m0_write         (ethernet_bridge_m0_write),         //      .write
		.m0_read          (ethernet_bridge_m0_read),          //      .read
		.m0_byteenable    (ethernet_bridge_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (ethernet_bridge_m0_debugaccess)    //      .debugaccess
	);

	ethernet_system_tse_mac tse_mac (
		.ff_tx_data  (sgdma_tx_out_data),                                               //                      transmit.data
		.ff_tx_eop   (sgdma_tx_out_endofpacket),                                        //                              .endofpacket
		.ff_tx_err   (sgdma_tx_out_error),                                              //                              .error
		.ff_tx_mod   (sgdma_tx_out_empty),                                              //                              .empty
		.ff_tx_rdy   (sgdma_tx_out_ready),                                              //                              .ready
		.ff_tx_sop   (sgdma_tx_out_startofpacket),                                      //                              .startofpacket
		.ff_tx_wren  (sgdma_tx_out_valid),                                              //                              .valid
		.ff_tx_clk   (ethernet_subsys_clk_in_clk),                                      //      receive_clock_connection.clk
		.ff_rx_data  (tse_mac_receive_data),                                            //                       receive.data
		.ff_rx_dval  (tse_mac_receive_valid),                                           //                              .valid
		.ff_rx_eop   (tse_mac_receive_endofpacket),                                     //                              .endofpacket
		.ff_rx_mod   (tse_mac_receive_empty),                                           //                              .empty
		.ff_rx_rdy   (tse_mac_receive_ready),                                           //                              .ready
		.ff_rx_sop   (tse_mac_receive_startofpacket),                                   //                              .startofpacket
		.rx_err      (tse_mac_receive_error),                                           //                              .error
		.ff_rx_clk   (ethernet_subsys_clk_in_clk),                                      //     transmit_clock_connection.clk
		.address     (tse_mac_control_port_translator_avalon_anti_slave_0_address),     //                  control_port.address
		.readdata    (tse_mac_control_port_translator_avalon_anti_slave_0_readdata),    //                              .readdata
		.read        (tse_mac_control_port_translator_avalon_anti_slave_0_read),        //                              .read
		.writedata   (tse_mac_control_port_translator_avalon_anti_slave_0_writedata),   //                              .writedata
		.write       (tse_mac_control_port_translator_avalon_anti_slave_0_write),       //                              .write
		.waitrequest (tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest), //                              .waitrequest
		.clk         (ethernet_subsys_clk_in_clk),                                      // control_port_clock_connection.clk
		.reset       (rst_controller_reset_out_reset),                                  //              reset_connection.reset
		.rgmii_in    (tse_conduit_connection_rgmii_in),                                 //            conduit_connection.export
		.rgmii_out   (tse_conduit_connection_rgmii_out),                                //                              .export
		.rx_control  (tse_conduit_connection_rx_control),                               //                              .export
		.tx_control  (tse_conduit_connection_tx_control),                               //                              .export
		.tx_clk      (tse_conduit_connection_tx_clk),                                   //                              .export
		.rx_clk      (tse_conduit_connection_rx_clk),                                   //                              .export
		.set_10      (tse_conduit_connection_set_10),                                   //                              .export
		.set_1000    (tse_conduit_connection_set_1000),                                 //                              .export
		.ena_10      (tse_conduit_connection_ena_10),                                   //                              .export
		.eth_mode    (tse_conduit_connection_eth_mode),                                 //                              .export
		.mdio_out    (tse_conduit_connection_mdio_out),                                 //                              .export
		.mdio_oen    (tse_conduit_connection_mdio_oen),                                 //                              .export
		.mdio_in     (tse_conduit_connection_mdio_in),                                  //                              .export
		.mdc         (tse_conduit_connection_mdc)                                       //                              .export
	);

	ethernet_system_sgdma_rx sgdma_rx (
		.clk                           (ethernet_subsys_clk_in_clk),                             //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),                        //            reset.reset_n
		.csr_chipselect                (sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (sgdma_rx_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (sgdma_rx_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (sgdma_rx_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (sgdma_rx_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (sgdma_rx_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (sgdma_rx_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (sgdma_rx_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_rx_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (sgdma_rx_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (sgdma_rx_csr_irq_irq),                                   //          csr_irq.irq
		.m_write_waitrequest           (sgdma_rx_m_write_waitrequest),                           //          m_write.waitrequest
		.m_write_address               (sgdma_rx_m_write_address),                               //                 .address
		.m_write_write                 (sgdma_rx_m_write_write),                                 //                 .write
		.m_write_writedata             (sgdma_rx_m_write_writedata),                             //                 .writedata
		.m_write_byteenable            (sgdma_rx_m_write_byteenable),                            //                 .byteenable
		.in_startofpacket              (tse_mac_receive_startofpacket),                          //               in.startofpacket
		.in_endofpacket                (tse_mac_receive_endofpacket),                            //                 .endofpacket
		.in_empty                      (tse_mac_receive_empty),                                  //                 .empty
		.in_data                       (tse_mac_receive_data),                                   //                 .data
		.in_valid                      (tse_mac_receive_valid),                                  //                 .valid
		.in_ready                      (tse_mac_receive_ready),                                  //                 .ready
		.in_error                      (tse_mac_receive_error)                                   //                 .error
	);

	ethernet_system_sgdma_tx sgdma_tx (
		.clk                           (ethernet_subsys_clk_in_clk),                             //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),                        //            reset.reset_n
		.csr_chipselect                (sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (sgdma_tx_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (sgdma_tx_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (sgdma_tx_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (sgdma_tx_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (sgdma_tx_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (sgdma_tx_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (sgdma_tx_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_tx_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (sgdma_tx_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (sgdma_tx_csr_irq_irq),                                   //          csr_irq.irq
		.m_read_readdata               (sgdma_tx_m_read_readdata),                               //           m_read.readdata
		.m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),                          //                 .readdatavalid
		.m_read_waitrequest            (sgdma_tx_m_read_waitrequest),                            //                 .waitrequest
		.m_read_address                (sgdma_tx_m_read_address),                                //                 .address
		.m_read_read                   (sgdma_tx_m_read_read),                                   //                 .read
		.out_data                      (sgdma_tx_out_data),                                      //              out.data
		.out_valid                     (sgdma_tx_out_valid),                                     //                 .valid
		.out_ready                     (sgdma_tx_out_ready),                                     //                 .ready
		.out_endofpacket               (sgdma_tx_out_endofpacket),                               //                 .endofpacket
		.out_startofpacket             (sgdma_tx_out_startofpacket),                             //                 .startofpacket
		.out_empty                     (sgdma_tx_out_empty),                                     //                 .empty
		.out_error                     (sgdma_tx_out_error)                                      //                 .error
	);

	ethernet_system_descriptor_memory descriptor_memory (
		.clk         (ethernet_subsys_clk_in_clk),                                     //   clk1.clk
		.address     (descriptor_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect  (descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken       (descriptor_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata    (descriptor_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write       (descriptor_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata   (descriptor_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable  (descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                                 // reset1.reset
		.address2    (descriptor_memory_s2_address),                                   //     s2.address
		.chipselect2 (descriptor_memory_s2_chipselect),                                //       .chipselect
		.clken2      (descriptor_memory_s2_clken),                                     //       .clken
		.readdata2   (descriptor_memory_s2_readdata),                                  //       .readdata
		.write2      (descriptor_memory_s2_write),                                     //       .write
		.writedata2  (descriptor_memory_s2_writedata),                                 //       .writedata
		.byteenable2 (descriptor_memory_s2_byteenable),                                //       .byteenable
		.clk2        (ethernet_subsys_clk_in_clk),                                     //   clk2.clk
		.reset2      (rst_controller_reset_out_reset)                                  // reset2.reset
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (11),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (11),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) ethernet_bridge_m0_translator (
		.clk                   (ethernet_subsys_clk_in_clk),                                            //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                     reset.reset
		.uav_address           (ethernet_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (ethernet_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (ethernet_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (ethernet_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (ethernet_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (ethernet_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (ethernet_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (ethernet_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (ethernet_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (ethernet_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (ethernet_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (ethernet_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (ethernet_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (ethernet_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (ethernet_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read               (ethernet_bridge_m0_read),                                               //                          .read
		.av_readdata           (ethernet_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (ethernet_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (ethernet_bridge_m0_write),                                              //                          .write
		.av_writedata          (ethernet_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (ethernet_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                  //               (terminated)
		.av_begintransfer      (1'b0),                                                                  //               (terminated)
		.av_chipselect         (1'b0),                                                                  //               (terminated)
		.av_lock               (1'b0),                                                                  //               (terminated)
		.uav_clken             (),                                                                      //               (terminated)
		.av_clken              (1'b1)                                                                   //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (11),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) tse_mac_control_port_translator (
		.clk                   (ethernet_subsys_clk_in_clk),                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (tse_mac_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (tse_mac_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (tse_mac_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (tse_mac_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (tse_mac_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (11),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sgdma_rx_csr_translator (
		.clk                   (ethernet_subsys_clk_in_clk),                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sgdma_rx_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sgdma_rx_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sgdma_rx_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sgdma_rx_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sgdma_rx_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (11),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sgdma_tx_csr_translator (
		.clk                   (ethernet_subsys_clk_in_clk),                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sgdma_tx_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sgdma_tx_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sgdma_tx_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sgdma_tx_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sgdma_tx_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_descriptor_read_translator (
		.clk                   (ethernet_subsys_clk_in_clk),                                                  //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_rx_descriptor_read_read),                                               //                          .read
		.av_readdata           (sgdma_rx_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_rx_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_descriptor_write_translator (
		.clk                   (ethernet_subsys_clk_in_clk),                                                   //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                     reset.reset
		.uav_address           (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write              (sgdma_rx_descriptor_write_write),                                              //                          .write
		.av_writedata          (sgdma_rx_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                         //               (terminated)
		.av_byteenable         (4'b1111),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_read               (1'b0),                                                                         //               (terminated)
		.av_readdata           (),                                                                             //               (terminated)
		.av_readdatavalid      (),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.av_debugaccess        (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_descriptor_read_translator (
		.clk                   (ethernet_subsys_clk_in_clk),                                                  //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_tx_descriptor_read_read),                                               //                          .read
		.av_readdata           (sgdma_tx_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_tx_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_descriptor_write_translator (
		.clk                   (ethernet_subsys_clk_in_clk),                                                   //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                     reset.reset
		.uav_address           (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write              (sgdma_tx_descriptor_write_write),                                              //                          .write
		.av_writedata          (sgdma_tx_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                         //               (terminated)
		.av_byteenable         (4'b1111),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_read               (1'b0),                                                                         //               (terminated)
		.av_readdata           (),                                                                             //               (terminated)
		.av_readdatavalid      (),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.av_debugaccess        (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) descriptor_memory_s1_translator (
		.clk                   (ethernet_subsys_clk_in_clk),                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (descriptor_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (descriptor_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (descriptor_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (descriptor_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (descriptor_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_BEGIN_BURST           (66),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.PKT_BURST_TYPE_H          (63),
		.PKT_BURST_TYPE_L          (62),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_TRANS_EXCLUSIVE       (52),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (70),
		.PKT_THREAD_ID_H           (72),
		.PKT_THREAD_ID_L           (72),
		.PKT_CACHE_H               (79),
		.PKT_CACHE_L               (76),
		.PKT_DATA_SIDEBAND_H       (65),
		.PKT_DATA_SIDEBAND_L       (65),
		.PKT_QOS_H                 (67),
		.PKT_QOS_L                 (67),
		.PKT_ADDR_SIDEBAND_H       (64),
		.PKT_ADDR_SIDEBAND_L       (64),
		.ST_DATA_W                 (82),
		.ST_CHANNEL_W              (3),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) ethernet_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk              (ethernet_subsys_clk_in_clk),                                                     //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.av_address       (ethernet_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (ethernet_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (ethernet_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (ethernet_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (ethernet_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (ethernet_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (ethernet_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (ethernet_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (ethernet_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (ethernet_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (ethernet_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                          //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                           //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                        //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                  //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                    //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                           //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) tse_mac_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (ethernet_subsys_clk_in_clk),                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                               //                .channel
		.rf_sink_ready           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ethernet_subsys_clk_in_clk),                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sgdma_rx_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (ethernet_subsys_clk_in_clk),                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                       //                .channel
		.rf_sink_ready           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ethernet_subsys_clk_in_clk),                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sgdma_tx_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (ethernet_subsys_clk_in_clk),                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src2_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_src2_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_src2_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_src2_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src2_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src2_channel),                                                       //                .channel
		.rf_sink_ready           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ethernet_subsys_clk_in_clk),                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk              (ethernet_subsys_clk_in_clk),                                                           //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_003_src0_valid),                                                        //        rp.valid
		.rp_data          (rsp_xbar_demux_003_src0_data),                                                         //          .data
		.rp_channel       (rsp_xbar_demux_003_src0_channel),                                                      //          .channel
		.rp_startofpacket (rsp_xbar_demux_003_src0_startofpacket),                                                //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),                                                  //          .endofpacket
		.rp_ready         (rsp_xbar_demux_003_src0_ready)                                                         //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk              (ethernet_subsys_clk_in_clk),                                                            //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.av_address       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_003_src1_valid),                                                         //        rp.valid
		.rp_data          (rsp_xbar_demux_003_src1_data),                                                          //          .data
		.rp_channel       (rsp_xbar_demux_003_src1_channel),                                                       //          .channel
		.rp_startofpacket (rsp_xbar_demux_003_src1_startofpacket),                                                 //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),                                                   //          .endofpacket
		.rp_ready         (rsp_xbar_demux_003_src1_ready)                                                          //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk              (ethernet_subsys_clk_in_clk),                                                           //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_003_src2_valid),                                                        //        rp.valid
		.rp_data          (rsp_xbar_demux_003_src2_data),                                                         //          .data
		.rp_channel       (rsp_xbar_demux_003_src2_channel),                                                      //          .channel
		.rp_startofpacket (rsp_xbar_demux_003_src2_startofpacket),                                                //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_003_src2_endofpacket),                                                  //          .endofpacket
		.rp_ready         (rsp_xbar_demux_003_src2_ready)                                                         //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk              (ethernet_subsys_clk_in_clk),                                                            //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.av_address       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_003_src3_valid),                                                         //        rp.valid
		.rp_data          (rsp_xbar_demux_003_src3_data),                                                          //          .data
		.rp_channel       (rsp_xbar_demux_003_src3_channel),                                                       //          .channel
		.rp_startofpacket (rsp_xbar_demux_003_src3_startofpacket),                                                 //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_003_src3_endofpacket),                                                   //          .endofpacket
		.rp_ready         (rsp_xbar_demux_003_src3_ready)                                                          //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) descriptor_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (ethernet_subsys_clk_in_clk),                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                              //                .channel
		.rf_sink_ready           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ethernet_subsys_clk_in_clk),                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	ethernet_system_addr_router addr_router (
		.sink_ready         (ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ethernet_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ethernet_subsys_clk_in_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_src_valid),                                                          //          .valid
		.src_data           (addr_router_src_data),                                                           //          .data
		.src_channel        (addr_router_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                     //          .endofpacket
	);

	ethernet_system_id_router id_router (
		.sink_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (ethernet_subsys_clk_in_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                             //       src.ready
		.src_valid          (id_router_src_valid),                                                             //          .valid
		.src_data           (id_router_src_data),                                                              //          .data
		.src_channel        (id_router_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                        //          .endofpacket
	);

	ethernet_system_id_router id_router_001 (
		.sink_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (ethernet_subsys_clk_in_clk),                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                 //       src.ready
		.src_valid          (id_router_001_src_valid),                                                 //          .valid
		.src_data           (id_router_001_src_data),                                                  //          .data
		.src_channel        (id_router_001_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                            //          .endofpacket
	);

	ethernet_system_id_router id_router_002 (
		.sink_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (ethernet_subsys_clk_in_clk),                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                 //       src.ready
		.src_valid          (id_router_002_src_valid),                                                 //          .valid
		.src_data           (id_router_002_src_data),                                                  //          .data
		.src_channel        (id_router_002_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                            //          .endofpacket
	);

	ethernet_system_addr_router_001 addr_router_001 (
		.sink_ready         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ethernet_subsys_clk_in_clk),                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	ethernet_system_addr_router_001 addr_router_002 (
		.sink_ready         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ethernet_subsys_clk_in_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                             //          .valid
		.src_data           (addr_router_002_src_data),                                                              //          .data
		.src_channel        (addr_router_002_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                        //          .endofpacket
	);

	ethernet_system_addr_router_001 addr_router_003 (
		.sink_ready         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ethernet_subsys_clk_in_clk),                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                            //          .valid
		.src_data           (addr_router_003_src_data),                                                             //          .data
		.src_channel        (addr_router_003_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                       //          .endofpacket
	);

	ethernet_system_addr_router_001 addr_router_004 (
		.sink_ready         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ethernet_subsys_clk_in_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                             //          .valid
		.src_data           (addr_router_004_src_data),                                                              //          .data
		.src_channel        (addr_router_004_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                        //          .endofpacket
	);

	ethernet_system_id_router_003 id_router_003 (
		.sink_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (ethernet_subsys_clk_in_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                         //       src.ready
		.src_valid          (id_router_003_src_valid),                                                         //          .valid
		.src_data           (id_router_003_src_data),                                                          //          .data
		.src_channel        (id_router_003_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                    //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (70),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (82),
		.ST_CHANNEL_W              (3),
		.VALID_WIDTH               (3),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (ethernet_subsys_clk_in_clk),     //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~ethernet_subsys_reset_in_reset_n), // reset_in0.reset
		.clk        (ethernet_subsys_clk_in_clk),        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_in1  (1'b0),                              // (terminated)
		.reset_in2  (1'b0),                              // (terminated)
		.reset_in3  (1'b0),                              // (terminated)
		.reset_in4  (1'b0),                              // (terminated)
		.reset_in5  (1'b0),                              // (terminated)
		.reset_in6  (1'b0),                              // (terminated)
		.reset_in7  (1'b0),                              // (terminated)
		.reset_in8  (1'b0),                              // (terminated)
		.reset_in9  (1'b0),                              // (terminated)
		.reset_in10 (1'b0),                              // (terminated)
		.reset_in11 (1'b0),                              // (terminated)
		.reset_in12 (1'b0),                              // (terminated)
		.reset_in13 (1'b0),                              // (terminated)
		.reset_in14 (1'b0),                              // (terminated)
		.reset_in15 (1'b0)                               // (terminated)
	);

	ethernet_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (ethernet_subsys_clk_in_clk),        //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //           .endofpacket
	);

	ethernet_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (ethernet_subsys_clk_in_clk),        //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	ethernet_system_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (ethernet_subsys_clk_in_clk),            //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	ethernet_system_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (ethernet_subsys_clk_in_clk),            //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	ethernet_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (ethernet_subsys_clk_in_clk),            //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	ethernet_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (ethernet_subsys_clk_in_clk),            //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	ethernet_system_cmd_xbar_demux_001 cmd_xbar_demux_002 (
		.clk                (ethernet_subsys_clk_in_clk),            //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	ethernet_system_cmd_xbar_demux_001 cmd_xbar_demux_003 (
		.clk                (ethernet_subsys_clk_in_clk),            //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	ethernet_system_cmd_xbar_demux_001 cmd_xbar_demux_004 (
		.clk                (ethernet_subsys_clk_in_clk),            //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	ethernet_system_cmd_xbar_mux_003 cmd_xbar_mux_003 (
		.clk                 (ethernet_subsys_clk_in_clk),            //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src0_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_004_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	ethernet_system_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (ethernet_subsys_clk_in_clk),            //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_003_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_003_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_003_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_003_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_003_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_003_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_003_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_003_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_003_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_003_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_003_src3_endofpacket)    //          .endofpacket
	);

endmodule
